module gw_gao_top(
    clk_50M_c,
    \led_c[3] ,
    \led_c[2] ,
    \led_c[1] ,
    \led_c[0] ,
    clk_50M,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input clk_50M_c;
input \led_c[3] ;
input \led_c[2] ;
input \led_c[1] ;
input \led_c[0] ;
input clk_50M;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire clk_50M_c;
wire \led_c[3] ;
wire \led_c[2] ;
wire \led_c[1] ;
wire \led_c[0] ;
wire clk_50M;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top u_ao_top(
    .control(control0[9:0]),
    .data_i({clk_50M_c,\led_c[3] ,\led_c[2] ,\led_c[1] ,\led_c[0] }),
    .clk_i(clk_50M)
);

endmodule
//
// Written by Synplify Pro 
// Product Version "N-2018.03G-Beta6"
// Program "Synplify Pro", Mapper "mapgw, Build 1086R"
// Mon Oct  8 09:41:35 2018
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\c:\gowin\1.8\synplifypro\lib\generic\gw1n.v "
// file 1 "\c:\gowin\1.8\synplifypro\lib\vlog\hypermods.v "
// file 2 "\c:\gowin\1.8\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\c:\gowin\1.8\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\c:\gowin\1.8\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\c:\gowin\1.8\ide\data\ipcores\gao_lite\gw_con\gw_con_parameter.v "
// file 6 "\c:\gowin\1.8\ide\data\ipcores\gao_lite\gw_con\gw_con_top_define.v "
// file 7 "\c:\gowin\1.8\ide\data\ipcores\gao_lite\gw_con\gw_con_top.v "
// file 8 "\c:\gowin\1.8\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
hpggv0Tm4wocDUFHdWKHHpAXB9LSbT6jwkjnxyWrCfCmz4QW6cwJlT3/UoeUCNUT5fJbIz9BfRVc
ncw6I5EDrnITof5tqjcfxkBgtB179czSfZnZ/ic9I+5tKSUSPz3yrZp2eFqR6maFJ4ZFO3ggJQRI
pMSxtGVtQNscosLDvlb7UBhCxLhz9HtSU3bAFqFdYJ6Ds4Gc6dUppvHj2vGY3kGoKWzRosBKS7op
WVhQl98MN1yzjocyiSTc23o5Z7CC4NoOElkZD+PHCv3QZatGCrF/Ixhyj7NkSJof9JAeqdxRN1Ol
uUZKkt8tieyz4Ng6dtNiWV1/w/P3xNM/Z9viyg==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
Wx+Z2F6166z7OXdCxTlURHlH51lrKlEw/V2tkTPJ4ddpwew0C7Mbi3RN/SMocOQTodX7RnpijzeW
Hrw2+8gA+9Mv3HskgEl+/CKPzSBbJO08rk5DbwzcxptXojpKt65aHNmSH3+/nZLR9U5OHJ7klLQs
X5gK5tvAHmk/f/dtB4WECVOVppFSFYyj8lGk4TRhh/t68x9Bwyu7SApWXSy7Y8cTXlRMfhDdDVp0
MjHTXirWWiYlRCUe43X3ZK6jYwQm9E5oXB4R1YevzbiMAhc5OMALYNVtBjnAr205F5RAnm2B8Zg7
T3KG+GLsMSyOxhOrJ01noNq7AIkMYL9q+hECGQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7072)
`pragma protect data_block
t84EYPKvQvKoQGITP5Is5fWsyOdSimIt8ClUYsC2dKvW3d5c20V/DUmb+BYtkPllhofqXOsJz3KA
Ke5d13ThaGEc2qPHxpE7jRDOimHBXF8t6BsaMFJFOsQPHT826bt4v/nqLr888n5F3bBw1Th29tPm
yKd+iA3Ob7qcXr+xKptJiyxGvxYb5fRlbIBAM8FR1yrV1ZrTpDXZnArEJDMQj3txVFUxl1PHSvwV
k7Ts0WSpM19qVLlAXaCpGndZzaPE+ncrpUcYBFvFBmiR+ULzwEJqEMqMZDEyeBXUvzpnQOJU+m2C
L5pDtDRXtbX/Wug/sNZG5/QfeXIjy4NbZxyOfFlO5Z6qvuQZSqlIAWcFcNwDAqR6/k3wxRoXhOUA
+EbJuNFYsXdn0TrQmeDlwSsVPRX3Bn06e4T+w5ZdYDfYLjZBFHQAZ6u5o6S7xhGm126u9NydoTUq
vCSIpicly1v4ONfYRCdQaNm57zBGV2oNs+GRp2PRprIPpQ1I08iH5Kjbzk/lE9VFFmB/Shjiawtm
703/XMbiq8wVJp5xMqrPLA1sj2GQx2Ijt30yF8xmS+0ZP/CkZ26w778Tz1XN4qJiFhP8jQckK5i4
DWRN+MrRM5jqrKQLec00dUIdYoRtQp9hrKufI1Ip2Nj5kd+WoHPA21EO47tZ3QTzW5+MEbcvy2XX
m/nISyub3fkbYzxebUyME9vCtO7+u6IOm47ty+w//gbRRm+hXY5vWdvGDLqI9+HBSzsYh4gt0Qe9
cOfXXw7Z/jPVdnJ/TFe9ffYpF0LDzmS7twlpESXx5pFhFtRJwZhz/00gepv1DpsdtGgUcC3YIhOh
ntb30QOgEwdTRSP+5waVEBj9M/WTj/6vSS6i9YtBQzwC7PlMabin+v4llg3SBQDplLCHZeo7hQXh
lTxAoOZeQkJBB8e9Zz3vHDaO6K832MKD3XjEj6OK8omnlBj3Q6ZXXlW6+EsfuFWX2yw5i919gUNi
qe/Cto5mJ3Ccst3OyWwrQzgMbPzzdH0U+KZGVNpx1S9mizaMSjLq5c9dxO34dmgYAhSdVJAK3ls5
JHyk7anhgHlmr0o8DG//PoJD/Fx+yBM1mWm03F7iXgqDxl0H+2MCosLRrCsYvy6Nole328lBdhwC
M9dm3orJue5sFI0niFacKkk1LECujmv3Tdb0jrtoK3IoXlZ2ZVTd10Fw7XjQVUXjZJDqk6hdZ5qA
s4dz0SbZ/O1KVq0COYD2/ufNLtxjQGF0OLeXB0TF3u1JeEJy6oeQXZB1i7R/MEwtXTiGF7fhM8I2
hHcqBOe70qFNFPMzb7f+l9U9hB7fdAooLkUXmnFNjbl3MfvApuNkAchbCS2Ec+SurDhTWXT/sc2h
+Zx5HxV6glQ5eMSScBt4wddARzUi+HNSzkY+8OqOegN/T3f3oLWA3UHle+LxJqawwz44WHXenK98
0wA++lwizt71U61Iny2wV9WYE5qn9WMY9yd+x9S7c4IrXWxcKQfxY3mpG49jUSYYyhxhYj7eWOFc
oIH8KvyJvC0hBJL1vOH7xOI48GY6RZGeVQZLIqapj10XYkPnpjS5/rITt/vPQkJjG0t12lchxu/W
NWaEouuLeVpywTPX/Gms7ATWLKY719siB/u8gyQhWfUTkh/TIvRrmFzbxUiDHzbdhHLCytw1WodX
Sjnn1Q601X1vqHFkEl5gWEM5rJPM2sKIRDsBJ7g3gakcDdBI/+3QOOHFxSSKJIFAlLw1+QyroFbS
+0nlITki1bzv5C0zjy+/G+iZ6oXwjG1BXhGn01uIrty00CobXlAPYyg5E8/ECa7QxgD5dbGUM2Do
pAH9/sbtVhlzAtlPDMyNjwTdnltaWeGrVHJ+JGyDw/Yc93KDXyKiInVm0vw6Olif92ESI9D9Ersr
w9wVtckRfzBvn6udsB/9OfVOnDaDWxwvnF7d+vhnDBhHoSFUc84JNEFYM1im/bpV1Rx4YDwsyQ6A
iBBuLXysTLXR4ggPqo+2fJk64ZDO0C6kjOHWb7zkKbOIWEnDI6mkagLKB/jRqMphY2z29G3oLtBm
f+KWXPKy4qnANnTw2qpKcQC+vPVBwlfqFtAgkW5HV29cMJ7a3EqaabiVTAuR2iU+9qJB9ucTjLzt
tvueaayQIiNwYkj6Xmu7ifmyBo4DeDnS9SCtAObpFbHFQzaVeksC7SEsCBl2yiKRblXabkCCyBcC
gXdfnp0Q2Lf4cAa/wrQGZGqfdIlFkgIgbZLVCU5KnXGflwDzq52e8LvUEr6ps4gWFP8QkDL1daSE
6wWjMJSlg9/RIF5UH4JvH/bVX++fJQXwNr7YKNNFbt9+nROIJK9H6FYRxPUGZMYVWmZhQd94XDQ8
NCsNkYi83mvhJgwj7DN+Zk3bs7bPOr2fWhI5HhmSnjHVKLe9LPkpS9z1bU5QQg8BT1QS9D4c0PuJ
oNsH4geoanPOjekiRaTgbgCjk6bRYnQFds9BOR3tWY3KPdmwM4bHNMpIxmtF/VtVO5UThi1gY5wz
aLftOHXiL6eoMsWs7LlgKNo/WvXDi8GyHT+/jfsScdUSojfoCPxp28rUOTgpx8G7AluOPP56eDaK
CtevhQSE6bn4OnViljHvarvS/3IsKMbd1XjIoBmkwxlYRltZrrlvr5FCC/+sHROwzgZfUvr1g/x7
yrdetspXhFl7fTiSKmHTKeNEd1ZuDKC+ZitN5Frv6mUyutkk+sJ0OBr8Br5BUkxkXyAv9avSokYH
3kde3O6x3u6QvU/1dFskRxA1mSl9XkxIy/7JwnbTudElbp7aeMMcQh2Lmn5P/tsoeXHmPrfaUR/T
PTjSJl+oOEWiynFNPyjR1yAJbg95/1AgV+Si+TkLJ2Kui6AXEkIQRqc/D/5AglaKLC8utp+nx4VW
Qh53Ln6ZCfhIw82wTDF/dOT/V5XAVnjes7EOKlpah0xPViJ3COZL4hJKRqrt/HT9F7SCOBGSf9hR
1ucMuaZovRNvUfxdts4myuwJAKuSUiaNv/089ocFqXO/T+7ZonJhoSpo1c9cbgpIwCxnLXUL6n1y
ZidwzRrBKslhrbAoXB0ErPLA0ObRWpP4N1H/jl188+ahUkbMiRRrZRoi4eE2yJ8tFeS7XX3i0tQJ
EMqTESeBJQIDVwrApx68ulA0FOMY8liC2KJm1LqQQ4ZNHUS4YBc5ZyGxWWRO00MesE8TbMdEKaRR
j9xyj5Y8JUdZlC/jKwTjf9Xd0B60g8ojZ7Fc3i3PltCmZxosb0spLM6pT7lFOk/RNY5la6b8Cize
xxJISuLngQRJBoedEl/FJtisCWSqlcFibOEUBwPJCRn5XWCCXMGnVmnT/qwTt8rwCegQUj4+noS7
PHpZLc81xjEkqm6G92seyYHcISOH9/zgz+0iDAJwwrI2dHJyIJfrnoht6dU5Vm87NI/UHdGUk1Gd
GYAOvVfJECaIbynJUA3itfd4PWjYHTF/6pdoUDcoctPjlloTM7ZEbDm/hCB6YZJsPSKCBmhEUThm
colmm1QDVMYe8PQNQaKXssoqG4s2XGkA0QLU9vZDJ7h06qbgIOdXI62Hvjyu+cfFC6vgAbkpYBhy
uKrXpiiST3OKuKRg58SSUWzTyQUG+6mf1CJe01gwdI7NU71HaBhPuieRq5YrJPFyDriznXsAdZtx
GnT6kuD77tAVt99EefIl1rNgZFmHKUYeAcAfMXCVaLWvwEZIOl3pHug3Otata92h7d5e5ZJ4sy4u
igcS9uMvCaVJ6LX58MjnOV5UPnYBCkMb0S2psKjjgSVlAQjfcDo1bvirgxPCUpILlc5CJcIl9/Rm
qEc6VGyckTtMFp/83dGoDffhhm+ij/AlgHisTkUPfEcvDXhGZBYC9gZZKI51YA2BO4d4C0OkzkKk
rlw0J9UQ68FjpudDTAJSuQq5EUVvZ5pn4K1215g3aNjC0Wq0x5yrhFGw80rbixV0bllQxXKsxPq+
/NUUFDghMectjl0ucJmJs72J+o6FFrUnEDW5YpFIoBhiLlSlSf/uKeiF4F+009a5bBxAJpIKah6L
o9eyIuptAMymQ2l7vqHqGGD2hBNhYGHYBB0ptgDJNOWzptC1vcj0pJvTQmCVujtfQHFw+kAnQWOQ
yZkkBWIRDxQNG71svR7EXQe/T91pU9JdgtXsCY7rpUV9cHKDPYyOo1M+qPCrSg0IHonbmiHFTiMK
VDKhb6LlvIuFf1kEDJYpTiZ31iGbxnPiEC+jfkJ/2uAzoXc5hiisL5eSCVdJoaWMEbdOrCjwC3b7
APTWPv5ChrJ6hPU0r6C/MGDIfvkG4emfsNuQIL/VJL2J+7fs0DHfWxc+b5mL69yI1+n1Y/lxEnh1
6B/IafrqKZD2VJp629a+pNqiFvV8KXubPv2Ufi/2NQ6qqXD9LF61aH+tjefwyIh4aYXcruuHIJrm
UotV6SYJZkVaHbUnjtoXgLACAzaOwoU3TkxcWAutVgeb9dseNabl7hNYdBdUROLWg4D7pNSsPK5C
d5J2aHM7+VEYd286PEwsIOI0IZuH+EEK/yQImani9hJtpwTTW5H3s9/ewmetkeurrpAD2BiSldW6
dUHQJd6BpZVvpy5TOgF4FogHHEeSnboOnoLbvOmSKpkSDB3zJETsRJf5xGn+omR1jjipko5hvNHn
znyu0TLs9j0giiWS0JQSs6FRPq98KRAVWETOC32CUKugRJMNlz1rMA2yq5RKJ7qvgs4dijC1reRH
tthNdf7++8+Wfc57UuCvgn+zFjbUroyFF4X7Alq6nC1ZjTOFc/K51lbsjVuLHf8406nk1zBLgCVd
g48h9MWCezGqhtfH/Y7jzLK/clKnc5B/1QSiZr54uq2FBuopi2dVVqWuFOeOQ+qR10A0eN5zIdVW
lbJbcks3vaYHozhiuFRz1eoKHK5Sy6thdmmNTB572P2qAeKZ9rPzWLlaRD2NiXIyGmYM1FlzvCzI
ytEi12Khf2J1+7+T1WhMShtdOPyM87+++ZoEpBQvoC7Cr8gIgPd3NOW7PwkgW+Zufjh1vkOLr2KR
kVLLxwTmZNnOiw8iaBoHoB667YgnTATemyS4O/c3bcXIqZ2vulISRRb2UbgTJTesyDfOiY9gwLGu
ynfbALUU7H183jqX7nGcQlWRiISvI8NMMwul6ct303PS58owHs93q0tIEaFT8kqlwLLdtZfpLCUU
L4cofyvAnDLV9R0woyLCAfeg2WGbh+25u4t9I7fKN65JB/pvWEZNpgslFdPfAkwU1WehUX35+ZsR
AXD0bm1FIZZzdkIHjvmk9WS+PCRaq3EcihGhp6HXU+0MX6UqhzlcCb87uivZpp4vctmXGwu6Z/0s
NV2z9rZ7eIgVluQ1MHWMNAKRrYMEbtIy6nHcbX5jBYn0y3RUrrhuMCZx2a3REbB/nXQFZQ7M18UW
5edvdQQZZ+B+IzSldaISu0Ufom5oCWXJoYxAawtUwTNOgnGHv7C2ITZ0eqkTle/LyaO6gz7fy0fe
wySZjMLzJ7Kg1iUdyCTuDl5n8xezy9p6R3kYiKlgoXXzeWsdcNmWXlzN0LqldhyP+A+eL9agbXVE
thOZPUmSj02vEndSkuPyswsj2R6Sf/Ov81TCQJd3SHfh5Evntl/zhRbN83WFCV3uOik0y+Vw9HO9
e51O/s+Jgv0cRn/3dDz5xN6KGGD0uS0Z3zfZhEdAyMFnFnQr0MVk163nP508vrbb3D8cBpb+BMHj
MtV1kjV6ty1z6KnhlODbSEJ1FN3kpBct8e2PSgUODa0YSo/bbqVL7hBGPt9Nxl/1S8HWpwA5hJmv
VG9x5eVB3kP4Hmol+2wXBKJJS3ZWL5Kryf3MXucuhRQP2P9ZFu2lGR6wMC5yuwONO5cpkSVTW1dN
jZQUO5RvBWlO7f7RSlBIXw6iXIc3LEji/HGPXscCpYx1I+jwzqhyBzw6y+1bogSxBwmeEDdvTMBZ
lCBhQwjEigomWSg/DZCHlGDWk94jXboOYXDrGdHw85NqC56emU5UiFi1viigF38QVARwy9zP3LV4
GaGlFQi12LeMjTYXuJbXAh29ziGvrYn5LA1P8oy2ZyLMK1AheF1PWMLm0k1ytSO+OKLFD2CIyQ4X
ncZmEQkKkqHQLRoV07MbX8GssVaViayrLiMQaDESer+7v7Ti5x78ti/ck2XmiPmAz49qZT3ugylq
ySmJThbklWy2kJzU/pIK26e3gb0649qrnV5Jjn6EKd8/ea1EUcDMxGBlNOi3AwNg4LrvrmNmrniX
mVh80r4EHCo7c/pvllLaY48SdcnukxuHctw5MoO48uJOZhzfxGtn1CK8gOiNqQmV2tzkcxhr5k/t
OXI6AVjWLUWtMfPc/eFvCC0yul76nKR9dRfRr3l0lUZCfiY2SqinP4XbLfzqm5nRAbSjan6vABZx
1wbarLUooUXCqgOc1agiKYlIvsXI0cuk7eKAxALIBP4tgD3mrSpB2FUj9bZGKw2BXoV5lDu+i3ok
4xlOaiMxc9k09gvILXrTcHeXT/wFHLqfld2M3bMoY/wJ1vSXILDCKq+k2EWowMT7DL0M6V7KtHpi
v2Psr7iCi3iWzNRv0D5TKflWtABOec3jXyCM6/Xth0Ts5lxq/d+biVb2Z552/bFrBoztamJ/EYp2
Y7Yx1mCxCvy3UjgpKfrV4gB4p7q22FlkGhX+z/YrraPolflvYthhNjWLjn55xFVVOe03hFdPKh9L
8Dsu5YqcRBbiyRwFQBmkXebfHZy7MGLgYthYuGn5gyjV1npCJwC3kz4PLqneYxSm0H60TjRpWyLz
uacxX06QhyITkCgMP7TGvp+r+71SP3hMSrQp5UmixBDhfO6Xt9d8zw+fryA9xUZyVroyhFa+JYs3
cKJjuyhNDd4bSllgKQpscmyvRp0+lt7FHfTZiI2WJjkmFCQ4yOIYFo1/phiXhgcX/U35cMYv+woh
b0JOm+1O4gqQzJ4LaTf6DqV1iWrfvQukg/SIR2Yoisq62o6qhb55DWLiDEQkJovEnBzsGxesSk6z
FlXpv6qtzpqOae9J2QtKv8mUAS7bPl73pk496uNnMfNsX5FFaA+WnjufX9JmFBjOxhvdVr8xd7kC
XNLFPo4+qh+9/NAYhAWVAAXVBWRmJ9SZrkc55M4uZ/wIuad2MkE8PtEPrdWCEZwmeTG+4l8OCwow
kNSA+Xa2kOBBfAudStqpCUaHuBtdiYKr8Ij1mwoqLxtWpHKzdoqSIf0s97/VcA8ZjkJtrZ63kcaU
WRo4KA72EO76tab5Cb3YSIysWZ90sNSSJrx7pVIixrMGavASf3CDD045KihM3eD/P6OZaxx9pJJW
6FModEbVfw8SGEtZl2OSv8ztBBrntCBvudThbWnw7t4nQRmNuQDidyj2dl/9tHSsiQ09JQtlInBR
b1OrFBISz0UVoyJOSN8+U28zA1t7dujDakIKT/r4FtEtICaEej6QwJxj0lWCEWBIdpv3lUvcp+oZ
t3Vnt7sU1Ad4JmMj16hbuArgLFGcKDZVq4EG0RDhJWUIwPL/ZvuJgXOOga2FdloX1X7acqBDdRlu
EG/AfkCDhTamhKVEXoGxND4uC5eAQGCb3dJHzQia3aVw609Jdn8w4z25bnjkEn6fc5VM4NCB8oTV
ZUAa7S53RW41v0+W56UIz9aSiAuLxyRzTN78ZbJfecQSsoGyrIOZPVISgaTWa3s44e1qsEV9qpYK
22CUPDr2h9P828qhSFXozjyeJ6SRxa4n0c3wD6vkeqwd8Be7T/a5LfPUkSNxmpr1eaApw2fGnq2p
R3AySgl1pkLBaCsbX2mVlMky/QEHzs6b7oLno8fO5zTTEBMRrZPwzolqcYxuLZlm5V6dTAprluso
up2BKRkkLfYnr57nDY/5TrpsJz6EyNREzKvWRWlM39Og89MSQgAqj5Wi5/NoIGeQUQibu1+XE/Pr
PLTlu4QUAEvgHlLlbL8hXz6OrCSGbz4F1joffEBgPxFJMYEybUKXzVnUxAfABd2gJsSaePIfmvlM
1mqsYCgi86z+JIS8+1wNu/1p6UietBnon1WuhUIlCXPRah517r/TTVdRJrFqLYsi/JxQtWum/R/F
/P6rBZe2GHsQjbEo/uLM6kKy9Ao3mvCQ8pDQTf+ZWn2290swDoUozUkGz2OgTL7fSmkgmfvJ/qtS
KfEr8wr2fpPSdPN7g+/fQIbNH4dUI0CJUuu617yNHi2FwEPxRuZ+oZq0AfRJ2ZcRV8ZvsSeEUT7f
33Oo427f4pMd/bfHfZnDEd2WVcdQ1C39FcDoh2y4OftcEa0TLoNK2y6p03XxO75IAV1ovtNTWRZk
TjbTuHMoGgdVkKSmUwfYKe4yd/nClyT7jtYXQOaRVUXAfCXIydzObs157NhEsJCHnt7ODdbPnXuV
1lmD1HWUzQtkhBsn/4NYUieFLaVrBlP5JLnQ35/lIuGty6OxRzrJt3teHRkc2ZoIvK3GtaSqtp00
41GUWcC5I1qMvjaKWL64FThM5H8/N3uNRqbt2X848X4sybJyNs2eZ8YY0q9qyyfEbkt0dmPqUN9N
HeOWk3gXutnYm+OQBkZ9+Fz2hTd+Te0e/Jxxo3Mbf1TGML1kivxBOjBpG5HgMjlSoWcAFkDH4zaj
CMQ6geIU92sC53nsPorEa0fJZg4gTldsUuuQZuaQ91jLvL4mmwAbdIc6dSdaZiCLgdwDfVQUsB9K
IjPUhzWr2dLBi5fYsLOjx6PLBs5uJAfN7CRYSyuB4hV6j9OmQF6DTfYxYaPBcNjFMpGpPN+Aze1L
svXG7cHkJGu8AuNFalBMuaadoGPnQWGm82McSQkjfCsNJnMhySKvKwtW3r1A+vO1P9N9oTuJwH0G
nOAaO6ghyAQASoImLHy02bLN+bbrKp1BofHr2myVaovGdlhwCpunemVxzaBS6NteLa61xdrfO0hr
hjYweLucjiEtdLnl2PziiW79ox1QBz2pNhLnFxZW2hRn8MTgrpUZ+vHhxZl/gNctRJrI//+gnpr7
9spd8vCmA+mMdSoW5K8RmcwSwiCV5ucX1BDXS8zVjPkKn/ZqFUX+AgVCN5vJZUB1JVIh/Tr5knFv
+kayhJ33mjPhDHywStQjKhav7d7M13BaNPGJu/4h4zJjx32BPI7dVddDZzYyBS3xRfrF+ELFsjnc
Q8qsJuATJyxbYXojJyFPxp6HrloxT1iOZHG5s6mWV1UdqzgS/jp/r/7Lgwr4T0XGk5JhU7bAp9R/
ASOlIHV6zm9MLhO+/2tx/Ckpc0rb1amn2S3hsp2N+J0ndlRJQsz3NoHEyznsQqO1LKZd9DpBHUN9
2C4uYbIaHwYEgF5mGObrMbXaOZtwRcs4MBnXQGRfs1I7E+1cfzbzF8pugzKRnh25u0eYYfiYs/8l
iL2kMO+rjD5WkAlyGAlsJmj3PvzSdgUZqpkwFzGF27fuFuZsRXVbaxbF9vcivehLgKCQS0g5Yfil
wDJgqQ==
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "N-2018.03G-Beta6"
// Program "Synplify Pro", Mapper "mapgw, Build 1086R"
// Mon Oct  8 09:41:48 2018
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\c:\gowin\1.8\synplifypro\lib\generic\gw1n.v "
// file 1 "\c:\gowin\1.8\synplifypro\lib\vlog\hypermods.v "
// file 2 "\c:\gowin\1.8\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\c:\gowin\1.8\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\c:\gowin\1.8\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\c:\gowin\gowin-blink\impl\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\c:\gowin\gowin-blink\impl\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\c:\gowin\1.8\ide\data\ipcores\gao_lite\gw_ao_0\gw_ao_define.v "
// file 8 "\c:\gowin\1.8\ide\data\ipcores\gao_lite\gw_ao_0\gw_ao_mem_ctrl.v "
// file 9 "\c:\gowin\1.8\ide\data\ipcores\gao_lite\gw_ao_0\gw_ao_top.v "
// file 10 "\c:\gowin\1.8\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
BZEV0Y+pfwZ1iLqHtdcSZjF3FQg29rYBhR1hszXZzyeum47USi6+n6n2T7XEJNBhOEs9nSCkgYqu
+A5maIFrm5WXyPh1crTQgMwbBahEf3caVqkg8iWHmTS67KyOD7t9F9SzWOHQmz0AS/hSPP8HzYAk
jblwhgb0dHHEos6ep2XjwTf96j4NueqRu5+G8OT2NS6ot33uhxehy+/Rb35XAa8PN80mAIhaqV+5
QsHfYCXedIfaA8P6RHYvPVca/KN2nw5a6OppzqQF7tlYKjsrYYr3zV31wyvrVe8zxfyltOlNtwyt
rOpdaacqNhHNZkKWAekMlcyBRRd+n/dPm2y8tQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
JxOrtW1OA4JdYRylW3xW4UPTwTcLiysN1up1jozKCvVKs/GFgnxIzWZwYaF9Zo0SPeT2nLN1iz/m
3VKW9Otn1BFU3sjeDRg+KFlMIaq5WVga0rpR/UR+L+YLBYYVThD/+Jb5rshGP8zBjwM8bVCzDtXq
84Y+Ibe4N9+ZAEkigcmx00FhcsKhG6wJap7rGnGOHugzX2hgTJGjH8FbrrdQ64xD/45siurCbVqF
8jZYHtw3CgbO2JQLl5u9m2rsV5E3DDBUgKG15HTVaQBLMe8CRJwIgSj6RlMyomxQd+r47DRGfsgh
0UjWV3DqlUf76mTKR65dO7E9nyiC313KnLgSpA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=10384)
`pragma protect data_block
zX5KxvYzeal/TnYhoQN89lWU91dFMnNxbc1WgQuZR8EbzszH2JOyfnBxLN1LQn0i6FHkVKsqb8v6
cMLzQikvlif2lklmydLAidAlNRLWN+wHwxMtypGfV1bUKWjlpjtgFj4XCHZJX4P5Nssuh0EXxlWN
czIA6gBLYQi92VRTZkBNFBPjx8oRWfP9mS5LeTJEYKPgRb39dzQmQKh2S64d3g93uPz7ue/ILDQw
TNJFNEo/qsk7bMnZa7JBQPTVLkdOAtAxI4OmIi9d6Pi6cB5hvN8mxNdnOZ4i8fCN5Zr4IzylPwsc
ZZ6ddwmBTxeDk7w1u7HM1d5n+2be5rjIbMtkDxi4zgkVTUwwzbkUfSjqjqvWeAXcVWKgDrJ5pq5B
BYFVPfPzIAx3qFcOPuCu0tCKASX8Tirg1qlQleCR6aTVA11KK5Oaq+wRiFFKFh7qAmkeAtpczI5a
oXanbwiE5uQzvChTmB40zstFThm/EMp3QaiA0w8v0kwwuWOHM2kH7Kl0EJWKPoAuPrPN2qcXSlSp
ueEVFc2ff4sKp0sVHFewZ4XFvFj616+eCs1TR/EzgsOvJsRSxBMgTTI74gsZdXNQ0lSZE3y3fOfJ
ARjCrXpk7sSLSAC7U/PcuX4/vwqfDPZYclr8hn91sKF3LJqFJ+00YImGHP5HaJJtj22+qUc/4+WR
AF6XGZMSnTlJZeIfx0MwpH7zWliZ0+D9bVz72/frpxfHMUs8dhxulggCSqFw5BsAly88Lul+Myie
fJYf5u8Ygz2KyNs0PLq6qmEocZsQFAIVUPuqzxFSgDO5fjKIKCE28oHT0Etg1VJ5dkVg8darHh2b
PPf2eMRH6Rgj7QUxhbZu8n8K8Hzanqu3T+fjzjbaVm0UIZfMFBC9bfdRQ0h8NCeBaw+LgrratqL8
P8GnIfzSzLKBumKLxXLFs2VzfnzYgklQbwKi5TmiNAwcAH3/cob1JjrsO2wSMvB8TlIwgZoIDaQ0
UwQm8kOEmwueVg1p5jkhvoLMTTmUgCvpsaCxrPx+8pCkTFYBTNTvyRnCNPFXrb6Dbo22G7ltmLLC
mWqQq3BDL3xK4KgeE9cVs93xWTDtr3sCcKpCs7+5/sFlzeKhCqbGXOUCy7OI2ZjvTK1c5DuFtthC
tUJQyOHGdPm1LXIBdwxtJkG9yognU8Pp6Y0QXlRDs4Th3QTcgwpQHzdaql3iFigwFV0rC69LrLq/
pHPlqGl+unTD53Nxm3EBr2GqhZX2RBa2txC7L2Hv29YdBzv6tM6EUHBCDIauy86zz91JiaywCEw3
uNs2wXYJpwn2pgYIQ031vtM67H86Fz0N1rnVwLWqGUrh5TZOux1TlipsaQiZMNb/+hB1db2muj1/
dtLsv63bLcxtkU48Cm/XnpZZZq17n3YcTY++OSOHwozC7++KIxGO0XP9Gy4ArruBPhDfXptJsoZi
ufAq1usFla4CGFU18PbqG9Ez9++Uv7Yq0xuNM0alXK3TjB0XaZUMd3Xn7Ib+6Ra1I89ZxYVwwdU6
MMDAgyR+6Zi5adgXRitCqOrAv+Ep0uHmshIlQr68/HRyLOClvvtHgGwAA/peujQwjOj4eaRU9iIN
B1vLdk47J9fCogrrlP0RSwksD37YTQGkCwNLZ4DqiwSbI7KgX0pp9nc7YPl8x0/pkqAMaFud4swj
n/UUcAwqx/+AZzRdQtS7MmaNAzXu9xSmUDFSeaNcpAIkVjWx/C8UMSDrfbKfH5tgPdYmF7rtWn+5
HzhYYRC2aSJTWUDVLqfVImGtgH1+Id3im0gUxkZavhyMZtV2Nb3Yh0xXeZJMojO4M2EOZ/9RIwbR
/x6URWdl4xLXlOiTCcd+DNWT73VGTkiZ3HXc//3BJ2UtThH+U0AkGJuxSwZ9DfVXUgEuV1YPVl8z
fsHd0zGN9wuFDZDNC2dDjqhQa1IQU2C7SRBoCLYDV4SEO/VyokmNrhrxDfeTk1B9WpGwxqC+4nP3
iS07Xa/n9pVKiA3Z3IGtdI1c2LGhLWzA4NuTdxF/zFrh3FxImHz3UxKPkg6EUxQadvZ50v2wb1Eh
ylEPDa6vgIkNOEladB5UVenbbPWB5EnYw+Q1FTAonrXbdbrcRKJ3MzgsfElcc4Bu8unzKeO+uOaY
pk/hs8689FcDN3OCRHgrhvQ7cQtlvbz4iTlIP5GEn+++xNcx1bvlbbufg5elwsjkTXFqy6Pzb3Q/
EQPaYVFQnWxbpdnLNhc0irSTjVMU1W4YX1wxnDotATGeDfwsA1lyA1iGc7v816ipAgrr8c3Ynf9u
EuHDPZXlc8upSSu1/W+2k4NQXyZeZC2aCVlv2QfLKwa99SJ6nH0Oa9PGeXETLi4Vvds59gSJTk1C
+1/ftPzjz2sj4UxQL5Vsem99q+6VJxg05lELS+n5HpuLiiQhWT60dU8J7AZPBqoCz1V3MFuqTG09
UKe7I35rZmm8DZHx5Evk4ieNt/mKOUA8pM+utBTEWDh6/p/d26XJ2JA/PM/Tz/2fTwVHp09FsyGn
upWQgkYmy9V9LFsarxgij665UwgHecN75SCzeqG0Qfn6yhuRqaev4wVIxWcfLE2rWX6vxsHmMqdN
Ox4U8rTMnyQF6KKficZRfH1tydvrY2SXJXb9o2uB9+/fNObixBw8f3Ya3GkP+w4HhUv8VBmsXJ9R
2TaPPfwkUiWgrdUpAiW8qoN4nnPWB7mW8uqoWEZu/JlG2OtSYPTjF+LHilRo3nxXIykoPSLdgQ5h
1FB/Y66lZrPMYwV1O7ADa9RPTxkBXEVtRCnA7s6ZdzLSRz4PN4NXeeKqHy3UeZxzpWSvpawWe76x
EYs+BEb3a66A6w0SWRjwFs83dzJBqitIsKu4jMWcmNRoan8+iBcSusnKaeMv2jIjjPqedD0p3wep
VWszKPGM1ArYXFeG/+yRPpbk5rD8GOmS25wOKxKfLurxDjnTmhPYhi2ld7PCmCt2YHCy3xtmhFvD
FO8kJfpA7ls+g3/WMXVFDwu9JSYkc2GWQpn6Kb80jSraGg9w11T0o7VpWDP4YVpE1EbTD4p4nEmz
oTl4DmR8Q2qcExGSiz8heVLVqXxKj0dEzFWUefL9XcH3gh1Cn/QI+EKWJosHnWneT3z1XYs3CwGa
glZM7/3oXiMBM4jtgUNajZtgZHUVC8gfxJuigdgrWWcGqlElo+lYAPb0VVhaaRRbe9/lrRO6Ouyq
7X00NDXm+EfdKXKevVjEJlMKSlRTzVeuSuYf82MQgek/fyKx8DfvTnxmffC+AeOkgGPBoXhoT55f
DBrrB5brOxQXiSMzYqJw89FZordZ8RvNZRvCgLN8hrY5cRu5GZC0dtqNEAAg+C6FD0oFjBPx35+m
cLYksNHPwRVrTk6/gOmgDfYAmXwr0lxHzjErsBvEjtuIkV68cRsyUA9xzBI3pRtphCi9Roa7l+lm
EeAByfi9MD8KR4rOr5c+JYpRLKPd16ZyGPG5Zy6nhJqhurFtHiYkvXFsWchDmJyyCirje3Ad7YZz
VwiQsTmLM6nPmv8W5dVrR3jbJbOSQWapHHJQl7iypg6ERikUeaHNCVwlgjxYpDJKEIImd/S7uhoY
ERJmqQdZEIlDu/OewpuUu7xGGvRDhcqiafzOoqhcp0wGkmOIJwiR7nTIJht4p0th1Mjn6hBgKc2k
5QjEQHeExWVH7erpcgF4IIPyLgonJYiR/L/nXtumduLSpDiFuv/D5GU1CcrfQ9k/EwPxF1JrMABK
Y6PdyjXMEYoj+xbzsHCff+bjcJgKmZr8MR7s/Bi33apRTO5E0BOU0GWvcSB9eGQl2s76AC9AuGFE
FTexnEKV6mp32eGKba/bA/FvgXxPBku9ta51hJ02nX2fIVsbbhtIzcrVUBAZ5JoWSylikqmZGouD
BFJYb9J1PpADvRwOwa/mmhiOEqTG0NP2yMU+WdyWcmQeZteRbEvSkVgh2vgYBwbbfR+cFhNBvKxv
v6RrA+XDPh48mm4X+kvzb6/xc2WQBoVyHtO7jEvfSHMMgcOvGq7LsUY692DgkO72+QOvGUIereLJ
TZ3rQfkG/aXC1Y5GSpHNUGSnjbRUtnTr/Sctdzr9R0+Dtf2kAyQzBCDRzVnezNmbgm1ZoGvlyyVM
YrxWHRQQofiKVtDuwCMoIhPiX6Qcfy4YKSPnTlL0reJZdziv/JQXVv1Yi6mqxUBrjiZspBwFiNbb
/QM8w3HYBqFudgwygqlx1gV3XRzdlVcoRpr6ut4YlI471PJFdb1YaiO6Pw14bY7iARdEz0Ff3XZW
bt1q7cVXrSnSX929gVkSGT8XeQg1V1gZQGc/uF4b9sWfEy7Vtl4F4ci80cZb+xzEQwXih6fY/bpT
N63GXDMmaBthzJ6BJ2uQzCwcvgQfhhoF0oCCb1urx/whw/OHEbzwGWdiclW23oDqzb/vxfI/0VvD
qUqkLHHQUYWSLLTCFQSgwULTbOfGby+2qPckMwKJLgp+19IOXmUq3OuR/UDKWnMgp4b4ZyQxiVxI
TvC2FbeM3A+jiCYXbaXP/kqBW3vKuJ1svE15ZVbPvZB+wwgO9s1eljeNK8TnpJIZKSBDUHDMexsC
kheN6fJauaOUbD61WKmW3cB/76514J7VJvW8cbCDDZIPkYsaEojPTSW1bcbezOrxJw8Bh2SDbGwA
Yrf8P1qe/bDfmqyZCjCF9/iic9BAJxrDPqCFREshN9NhrDPdNv4t6IUXXz8CAzmnwQp8oftvgcQF
c99XzQeIDhSpLDzLpHCWCTYKI/I6rQ1JsVG3xgu8OQbS/puU4er4TccPGEB4j9tn5Xi34n3ncN4t
YU45mAtqmOlWNJwmK5PTaFbNAI//15+nJ69VtYKS0rllB16x2ogcQsjPCXEEemT07W8Yn9ra8c5x
p++yLNWm9DKg02cX6+MRke8max8CDtZ/PbS7JANSFvPnEjX3OFlfR7EGMOVTVSiorq6WDgrJNYrf
i3ON0Syj9ARbYRi78IrO4XwAu+TB0ehFazPKjplZrsB42PyL1a0rkFiGQ0Vk4i2rMUpqBHTfVqiK
ZHqsnPoiWFfjGbRaGEE4igK3mZOiQk4gXEJViO9hAXkFBVQkfM3njgJtIixZhG9QfF+QeQOWmJru
qZISml/p7lssiEd9Ys6KLAdxz7dDGJCVQPIBNJ5D/eOyNWql92t9xax/bOYoFLWLSNQqq90nsU2c
U2fdXH7G8Ui1/brIkrR2Qo+y8w1HyCM7z+L5Lc795G5225D7S7NiR7FVZWNRxYsox89iMjnhoPF0
b0ReAghEopr1HS4oM2/prVVCSuB8UVC2Q1p9Z/fXEo70ye28Sx8Vy80uUNZWuDtSCVH2AUpTHMxp
kzuw42i2Sq3g4nIW2Lkl8B83BmYYKRQGUJW1d+zK5I5n8Pz2K+jVorEk7qZJYGOt7ZWMlZVSHb+G
qkxpp1Ivl6sL9iXIAA47zMeSw7bW4cQAVdKVZBhKsrymP0J7jphTMUdRYfJJMGog9/iF0571p1nW
pzrFSIviv8DIJHI0nDXGEINpBr8kWrnzRvNFbflAh6wHOgY1PIkgOC/+mjju+0Opi6njZrxd9HEn
EdiDDySIE29JHMfmSpdsKAewuVDu0th1jAuR+e7VqiJ627jUGomFj/3QVcIoyoHmTQnGyEaMb+5y
XwGRtD4sbkiX87Sb0BeZQhQ/tgjo1qIWhgftxRXProw3k9Q0TJhd8xyi9pV/p33+F+8Cc6RqFBlA
pdVGKRZp2nTAUbzICZLYMAWmteE0xBQXUJ/4+M2saVs5vosKBvUgtMoO5Ock2904mjDgIdEHL0G1
QOiip/z7IpwveDd9GNdbVE3kJDUF5vEcY6046CtfPxts8UQqgwwZMTuG9Mx614ew2T4tDJo+UBst
g6d4dcEU1dGMdtCT800jL6875NHC/jxZgDsxQa7rlzSQdhEmjgTBWf2qj8K56FzFnx5EE4fgnY1E
rX+puEx1S9lAUV1vcwM9XgynOHrlnnrHLA1WWH4Mo5KjXpkTQb76nyeZhDC6VujvQIf3WA+4r7nj
0oCBucdhmE40v3hPcvUkrtBHlWG2SSp5i3hmAAFFCtaQ/EO9mKcYlvj/wRWXkApCm5M4rIEvmz+F
9kLzEpWe0kf8JEqbXK31uDF9phmDq0ja03xBisq66y2MDodQKdbWWraAcedtm48M+IOzPU9Y26kc
KNJrL3cr42uvfwKxGiCXYlzjSpPOucOUxbYZZQm/kCoKbTT+JshMe6TVAQJJIrx/oOCRHcH7uIr/
aYGQzI4pqEGZn9SrxzpvDbz5n3IE4zwtEeyIZmZ3lm9p0F4dXHFhpbPgMt7p1mmVuRBnXMWGsIqX
F2S3yEvf+6b7m4QSG8ec5qazNhuUfshPPF7EKK07i+N6YWm4DRpzeSCk2TMDteWAOXb8xYrH0+qq
fVQqakyr2NINc4kGtV0CyggyBWWpLBM6KgyLEf9g5xligHS+7lh9MshWg66Ij25EJ9xk2DwTrvHi
EVN7kE4PDzpH2mmcVeFcQH4NDOTyzhG9ctA352BH7wktwLiCXlqqNZdsUo4PLoKiBu/jEY41s+iW
5B+EaA1gFAqXnXsOEmAYjkWbQWP2XbB0ok7jaJmiGFLZD6cmVkg0wEpSX3NK1XSae2gY/+P+M6n0
jyIFqEGNFx6CPV0huyEyRIoFYBOOlhk8awjdXsxo8iGSAk1r6ryZISx786pLsPQg0EzBGIldOzXS
Ois9uZwX3hcQAeDzu9QxlguQHst4wjq1eiWYUmD/qbzbNqQzW4QPZi0JvGD0FjJ5uyfCRTZefNld
eOipf4Hp8l4Lh1DyJ6xCHK97L4UHZlJq+d4bou8Qxs+6l0XVgwjKgiP7xgsZEIZv1NohtS+0Pk6k
ybk+p2yuA1dPnWlB0fxq0FCi/Xa1eYSMYX/OdsVi9cBPDwfKtk0ivIrcKagyoIz+UMWHSKd4nqXK
LmXFxznBOPMMiKw0+Hp3R2y5vEJfjjyOPPrRzw3VqtTKdy5nIfGnYGHoeNPqsR7ciKBE+jx7zgKs
H6vPwHoteUp6fPF5+k3q0X5wuQ0eXgzetqgNGeRK6s/mCeVedLvOFNRWvpX/udGrQpRNyfAwbSFc
UrhfNCUBuZ7j+aACHl3aNVPnS8hv5rPTrPK8pgJUBmyZ7zFijiTsU9RWfoDW2xKmjTdljXSC5LEj
RHbLdSmjSnqrRx+nA1ze3GNWqjfAjxwOPxX0PfnTSaBaQfwbj/cMlHBs3KJZ/5tcRg56DTa/wnB/
HQapV6SVxedSlJe4lZn0b97vSWCt6rCrFdoGs++pl2LwPCeq0e7QF6iCBnfZAhO/lkWgwVCUnqHD
KrOA9b2RwVnPsaZUdbTho7ceu+mUFpr+Kup+dp8ZC5F3foAVToL9YDwispCwlZYMBMcisU7uY0YQ
qb6Klq9drxTAFBgsWJI0DLEXClHBn9cBSS6+M4Yrc0BkDheR75sbRm1fssubBFmK1YFS6UJvWTOH
uV+xI3sZmW4jrmzxgaUZQFhURV8z8DXC//EDS9z7ggQ8UE6s5bI0g8QukTKBGIV68hujkTLLiF5p
rPW3WYjI8bsCWMSgcPy6DGBq+wp0/anKQrX/IPXSgXcUoCOdqRFc5SxzDMdF2t2IXrCaaa/2KDN3
z6fQ+U8DALL0vbcCNnHIL3avnmFcnrAZ2ggNytVwgWdnov3VcWCBv9JtubsrN+vs7bXDDinGlOMD
D4+z9Tw45XJwC+SUDb7uO4Ki5ykmiAYx+HIvnBjgjwIDnHqMo+TGAVC5ySpRUB1PXa8ddC6f1zwc
2b7a+8EHK3CswpVc+rqzs2RYyXJ6QihzUFogc5SOMMuwkBOgbHS3fH5zZ/fHhU8nCXiaGEqcncIZ
+yqKmChMucYoI6lxzNcok5MaF38Pko3Dh5vRDahC7PgRc4SeZ0TZHIn9lpgIg8wDA+O7jiE+BpGg
AiZ2uqGU66nIQRZFVwTIFU80ihpb8ciPF4hzjBg7mtQpC4cZpNqPxY2O+E8/NBOm7D/tvWKIovT6
+6wbb1ZKa32G+lqJiSZtL4m/Sa3j/Phqi7rkICV0TuoLZ+UA44mcfrfEtpsmi2R5G6Ypw3pzUYXa
T+6QKnzJdjNHkzxjGUB4/t7H5VYoaylRigAGjYKkP7T0kdwMjDhV9ryxtdkogRtfbTcMh0d0rOvH
UhUGUI+1dpcGQvJD90qvJhmZYssFakalrFzRE+a6H6oZDxcJlvRpgDGxFNNP6UeWQ551CXhv61Ud
dEGU2DCVKlZU3Zth9MtHjmWgw9/WpLCtvC3+JhCuAQ5uEe8qUqKePTjEsnf7PXXPxKGJ0SuQMAGq
7mW13a9t8xwU1ADeW6w4onihAeF+sZeWPBNtmXei3TxTWxLjbstJhsrD87ug4vnPvoom2XlcR2Tl
SBO8Bi3QV+nCGbgMRMFmuX4kIo3M8rbW1sH56MnisE3mXR+fR9W2+tyCwwr9h553Ydcpi94H60HY
lnYP2ZNaOwJ60zpQ9DKkg5pbEAUJwubWlL3j2zCtxW3O+zekqX7ZEuydKbLjvQl9rtZRw1aApM+m
8QWGtKfbJkNK7tVyYcbmCJE6jJfApoz/02XtBf57s44l/bQ5qhfSv6pNb/NapRjph/JKamlh9X3D
yZzhXbF8T94WGKA7/NOXfVfUqvkrg+mrmEx5IicPmmnkjDsRLav3pzldxwVm8F0+pmQ0x8Gatl/2
lFgPwMwV+MBLvh1+3xXYWX0/i8UNXf+J+FhKBzMQGlhsjNbXj8yf8fyvdqk2n+7FKDBb9vbwiSOE
vYQBp6JugRDArQi7JPsRgxY7n7MgxrmYDJgZoCcJ/6tWSjWvoxx312GHE/u/u0SmgiLI4W1lj+ld
O0H5GYeLmBSWGFyNczqA0ISrtRdg1he2H4wMYiS5DBlrg6nPuGDhD1XhVPFE7oxLJZD9MxyHBHt9
YgX0LFbdyy+lnKW4FTQg4Uufg7Vk/iiv2H9xxoULlydIHrBN3RmstOFUGEaJxiycu/z5nkqwO2xK
7+ebA0HEJ4UUeUmD5dFEQa+EImQ5pufqwz+h+TAIlp8Zc0QnvaIYLi/ro7VYamwvBDFmowIggkIh
5t6lvALA5hhtb0IFQ2YDg2qw+ZfhKqGQDBiML5VZcXFLTW5Mhq8Qn+HkrayyYQqKlvRpxF29DEXx
exo6XDOlCVQbTxum18bpihCBbGS68zGnHTDHPSI4+tHLkHwxuztAAxNbob6W3tG4qg2/vI3mjDP8
tHzlt1aWbvQeOy85s38D49ufgU8agdXyUogsjS8JVBIj/I6iMHp0/By+wGg5pPy7DOiNHDx0UFYO
wq3lPgn/N4kR719j3VOAO46/iGn0lA7tms4UqjFE2WqWiebuCbLDXK1ktDxIEv+t7ppgah04P07K
yuv+vsdlvFqxPVAkgaVKPntXMSZVUsqgJHxrWmhz19Ang8rhhRTBY3CgFL/1mzKd6QP9FOScQhbt
FhxJYr/vDCAIl43JQ5of4uIkJu8ZAmguEPmlYipXyPeBQdQuugqNeVufLUkXVH4l1qa342zEldOK
4bPfzuqhKKV/ZQWk/VQCuefs0jZXrB4G5rtZK6E4mN3IAUWw3TQOK1JswjG/KiFGD2cCgV/lI+m3
DUVjmSSDme/ZIYjSbOW91oj4xmzSeX28TIaxoITabZLl0s3vUp8Hgyd0bGecWv8fUitQZWxYJxct
M6aPpq1d4FFHXMOfaqFONtc3WpyP4CkH7PtnbYPQ1ifGPtYOfY/6Huc9LzLCzvrrB4fnfLVtwRtw
pbS+ROkF7bAZ3ZDh0sHEEKF3Mhy8I0pAQIPsP8+bD+7Ddn6vIBl7xaX8vHyvbc4JxmAQELRu1g1t
R1gxgCR51/GeEdc4pzkdarlbWqCyTpGcojYIK94wn6emK8XMDG1FUid0Vv2XqgPQvUuo4pHN91Pr
W3i1/2wEqiuGWznXvEbiwZx3XNC54KsQe3TApQXBtLieV7nMwO6+2/cvDO4ZGjYRu5gVeWogMtfI
ssilbIr4doQUvd1xzBmrv3L5YirlhbiaambxnrQrAZATjqywkyLVydn6juYeJzRkrP4EN/vTowfA
fCV632H6N0DiFaNvphSjsLHAEyJqE+9p7YAg9zx66rxJWT2VmBZlp3cCDA3UijZaBPW6VZBnG150
N4SFqTHYTfqGMqQ3WU3AVG7a44yiQE/XMoimYaLjs/eebpXI8SFfmGnHGET38ObRVownP3T3Xacx
lncDYWe5CEMcM+n56LLSFkLuGpMrq+x8lmignhxC84c6XyQOA58qFX3Xomc2dUx1roU9oJtk3z8s
k/3VuwzZohO0N5KAAHw6KaqZG6OrjXh4c7V1N0WgiTej3XaCZXPBzu+MhQreWWUIBay/Q8M9DhgF
KY4gvzyvAp8tl/+r8MZuwSpf2Rx/zwGM1PypdQcaS+kAZx/ObmXQLmsk+WkQFOK0wfhbs5jTFcur
R6caeyJgc7QxbWyJqsqYWDncI4UKcVWmFP3az9xenv1EzdTF36TBcpN5p4DvMCHju8382JMAGyzP
fb9rmjJflwgOle1lMkbGNSp4KjVjxKw8AlWda+Jfmn6VItgtSf4WOPVSTvFofYuaJnGy4EPwEKFN
ZHXePvjz55o86KVX6sbEvIUm+vYiaYwVhgLRgu5jfelS2GZCLNY/d24UCBAdu3i6WviYF+ZmFXkc
VD1ZEUSI53E2Y5fOM/arS0sxFwoj3kXgQQ4qYiGT2ZF995ivym7tGHYDanx8M5xJcucvrJUYRcmr
3Kf61OuTVYXruQj3QJ7nNAbUsZbDDtCcnZh+i6Gtx5YobXYGcfahV9ykwWxqdTgdZN7XofHJ1PqH
1TYnBwSy5q+BNeaoqLYQ4k7hHYVxpKtC8jvMt0iMnmqogRFfRjHeF7Rlj/hGcA46+1oP2woTEzBp
VBVwqPspBnoJ6Fd4CuFNIAziwdwVk+tyMTcln82CQQ7hBMzbIlcMq90D0iXpiJr+DD0k976W5b70
nVW05okwNL8tOgpYma6ZJ48bhNnF8N2Wr5TVFoqXvx8dB0Kwrh/8Wsyxn7gXYe5jmHde3ZRJGfRn
6/ktYyOFQKTdalMFlAtDzMiump66pkcKC1u5WuIYXOBi7/SYY15qaKCnmGAejyLzSioDHbrxyzrz
hFEXVzZtOApEzT2bFoCFxIRhQo/OCjkC4img8G6QdXh5bB6JHw661tKpYtFTOF1NnsUqmCeMx401
H/Pxc4WKGdTJZOuvjihtEsSMnIglJWS/Q+hXe/n0NXxMWp3sx4vnaOkENda3w+y3H8Mgs3AqV9l9
uvIyzzEtRhinRfzoHxE/wK040g7Atv1xtiOc6em1RObIE356hIQb2GOVgPNlQZ68vlW5woUa499m
tiGJtAYcrYWtrbQ6cRiezmIelvCVg1bT7C9qZoKRZMK04WEkbQQOCa91ulW7w0ZSELbFeshEadwp
sroUa/a6WsLAFdPLGD2FmfE8Xcn8bEsjmk6EscWMzgLSMdRwdJixLMeq0DrpmgKyW6W21XycTOv5
GdHiaIUuMNkfXmw2WXDeLdPRTohd17W9w0E59JYnMb8jFOmSbcq6lbk/OkasjgzcXZ/737am9/DP
tN66xvBRbpBY5Tcx9J+oo8drdYdoZqxM8udYY1Hjdlk1Xe549NL18Q+LczP0KaDRofXJSqtMgjv6
Bw3ljm/Al4HqycqUIaZgagT1cPClm7IkPqhWecWgjPqEqrvoETznOUDxUwby04rPpn9s0LKu7YDK
RPjTWRSm0kMdAqhe5ncK3Fx6WXGmQDUNPsmJUFi49cqLwWAmplNjN+jEzcQSQ81xevhDs+m1MxyO
6bMZcMxbNtxDNrw1GMs1OwqKURL9fC1Hl8QI/8YxvHXNOv/LXSD1MZfpW+TS/G+WK75i3U2u/3Ak
K5tv23HH0RaqYwQulVhxiqPhi54D8G1BVghrb7ZrC7a5SiQefVprCiBxaxekF6IM9AOsaQ0V1ybb
zNcsbdKYbQ3H5yWgnNrtcDmctLrQwutQ+69Keo1jiNu7goCEL0xnJhWIQHUWmu2hZSDUTAJM82U5
dL4LfBzeijrxy1cAQcnb/K8eWHJh52t3TLEWU5X/P/83FHvD/JePkgTrVR+utd0GyNI7OiZBF/AQ
3NX9EBkyXhqMBy11pffSeU1QML7+Ae9ijqsfTi2RoTmG7O5jgnVyG7hgscyocWOnsnq7cQJpAP6k
qMzyi/mof9LPMYo74nYnt2KNMS8PR9wvOjHJ4b+ij4UGTS8YAOaKqlpK+fYhH9J9HgNgGGoDVJ0e
TAhYDIXbrFgB6Vh79a74ZGfFxD5jcMcIiB7+F9HOjbIlrtHC6NBxAfEt58znsjfEeDdhWnDFi13V
EBdazMPsGNl4HiZrZHswxFXMnIHiD/VLg9SVnatwT/D4YQIXqz3QtyyRIAmiCRNHpVMamJsAILIA
Tn0e4SxOv8xwLg9Vz7fDVPLKgfDT3pXoOI3/AaHzVO967VGVGSJHwL5HuZijFAFbHu9rmCE39m2A
gr8qKJO2vRCUoSZV5wwS7I553czXKNIcJSFAsL//gCcJnblIUNoHTgq/ztDkO3JylJpvHW5vlmBi
DLZ9iP7EDCiz9XFv0Enxi4a9W2Awo1oOq+qKTtwHvAZqXaWhpVMpuefjjezrHZ5O6eoy5Rvf8N+U
XUMQ8kqw2pYUdJBv4fBAWVtq7JoAIKNUsEU6LjeZM7F6Q24X/5l25G/yQUz/s4IqftE7bEzfmuSY
vg1viI/pxP5CJUqOrIzqnpYZun2Crz36Ot4x5PC6WOjR0shMo8glGAu1XfYjON/FvRcvthOugPrA
v5Gb77AMpkcpz7hC+1CkAzgpTbirKr0F95iiF0L8nF4cOhaHCMeee+yD3KQMMEvWBCGzpRSeLeh9
zX4x2R3/6sJP980xYE4XTZtUPGawtFqyOIL8DMl/vo1PjTtbNFew7YEOEqK8MLPCCxhudqlj1qeL
IUA7MU/LN4hSfhPWlVnLSHyXsqA5wKnwARHh8nSUlAxaUI2ZWqmJQIhJzV/1VG1K0tQjysgIu4sM
JsDVC6/qFlVTvdaHOFQlnf6ydZ/vVPxbYSLYw4MOXj+BuMipsLgrmVZZkBbpT98eNFTTJ4gIeu0x
4mBfunSKSRslSysVuKwyR054iI2CmHrGEwlJFB0UN72nJmoM+ePKay2AoepiY8uaPk1kX7+Sh+iG
JjP7pIJhoIAUg1wlGXqNmyzDmXrv/QpSUU1xVVQ5kZYwZIZ5x3yu11756lU3+kifoXTC6m7KTx02
EGUnia+EVgKh6eRyMOIds/5lxbCChnHgP0CiEmUDnqZGv9QWDwyqCRzgBRxz2BZ7ZS9ttLSCAl+l
3FAxdD6Kzj0KBTW2nkwcZIaW85DDv7645oqoaYBm7e1vu0E18dW2zDIfs7qECr2ljxF6jEXyapW3
zxX3Nb18/UZp9VZcbBmj6HVbS+r2+Wx1PojpBwyyAHDQWK/uvx96MrHsehaw55nnZiyGz1xRkfh4
ERidKbe0Bj0bHbuqLN3GnXxSYx0fgJkQ0LWJJE1rTb4rljoynzcv4YjBFELaZY2MTRo8pILdLl3a
d49G/MJ7rAIpKj3ZYBEMmFhnTFF4qYpcvpO7Ai+SQdntAXSMk9TeZ9A0SJf2NxIeT5lNx+x6+aeO
w8G3InGIqJ1BNpcPuwbalMxZkk7JFxFq6E4GqxaoudhK5UEnu3RF8faotK464t58X6l/QXXHnszH
r/rISSkw9+f2/TP/lLi4LOj1lriPW36pl/zeUqC53L4AfsfJM9vmVevXXqw22gVyBSvDK8mqqPt6
MsuO2cZzEOxLBSBpunvb2Gz+1hj4TcQlv8wqk/lDJFnbnoTST5wyeU4HrkFxFqSVM7YwW6uTv8LM
O6ZyibEwjBEjiA==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Pyc+7kvzBVq4Dd1VwzRmVBEktK4e9BkxAwVgiiMBP4OI1yNwt7F+yQEhFvLcVH5FBU9k3Bk5g0R/
fGNscjfC54DAtJYGJoHSC2Qkju273ZDGQ5GBZeBA+Omz0LR4NGnYlrPzdj7g+x/czmcW4gPDkSLi
1d6y/BDFhoCYzVB9BJYMvhU2yyBd8pSDDskw7+4pB++GO3YMxSMQnAsSP4H11ROUUPSYWSz7Istd
JaaSkZFuL/Y+3gs/NCzDvX+aH2rt7FrsNAycbWtUKp/uPnA2vMEBHW1/ptnWFCfJFCvStvn4NF2b
o+bFlc/NfBYrCvp3l8g9z22fvrCKnVbJ66MTQw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
eIBgxZG6vpy8I9T7tgjyHHEL2Oagvj/TL61YE18ebOJrz/ONyRnM5TlDVcd4ieAcUgFStMRfiQAG
9PK7xF+45XZqhdWGzqcb8jHcqb3sqCjw9DKlKwnGSZfjC2sYwUpwY1a0sIEPJHcJKqWdB9fXqYAu
p0IEwvUF+FEivmc/v5dZQFWtUkkXSXNRuhbEGrFbKFeRoN069X7Pu7Q7ZekQinv0IeG4PTyASoE2
KGB5b5bTQeuJWkqjG5PorXwKnmAQiDQPvYmu1gBHXarwUU4flYl7hQnm+THGy5clL54o5zDTb/m+
cY477QNFS3rATN3G7wlvwku7f2ZhcCBbeXoJjg==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=58960)
`pragma protect data_block
9sPS9Ov16O9vLdpiDrePMvQWxnqG5a4tiEdF9Hcyfcqi/DJdXZJWLuUV9SbR9Iiei9XucC83wyxM
+1dlzYFBrNTwFVC9QMKTGVKX6wYPIYczxODaUVESl5i0FTR8Xgud/VYYZk77XwxURxVVTAsSJ3U3
lVuYWSoIPYJ68iew9+DgPxtCLYFySpV6EeLNmBeUah0bl4bnSm8DSICeZeAcJE1jNQUE9m/94ZTH
Qos4DbNdzWZyaD754QrcURE99qTjpzpiRISoNl6b19+gguiqpnFaMakJzmHLTIvqQ9F2f0NHVgtE
EVfr1yqJ4Pgk9owqYZBlrlYNQbdy6lu4wBdAbFlIjxdQGUy4zLh9+WmAV8EarraT7E2IAADbTJ2v
cNWhiBVUGmCDm9kgi7/Z1A0k4mv/Iqi/IZHedCidabTfFhupRVVdZMIOM3K0WpDUqJvdPcwax3YO
WGtzRVEaVdMo+YixbY3RgjnDe5uOC7tEYNF9kBa46p8yAmHjLlpE3OTAoqEwyd0TInd01kyRxU5q
oZQaCp6ux1y9810LWOh2Q5wxq1WuyKthv1tpCXdP7HUz0qayXlJelDRb+zB08J3GaDTPMF6mK13t
kpSDx2rhgC5IF+gQEQeb3+pyXS75zCDW5LYbMD12Z9aMbwjeGQeyuXuBS8BqexUD4Ry7eA/NMvzx
QnsrA8I0YrX6X245iRn4AkwDtXkGuI+IgLlPRjPE/VehFjOodBnlOpCmq84JsCZMpwoACcgfblOx
DQg1lGyLoe2Qnvh0YRRUvtHrapN8hImdcG1D9hm9r4ANiKkAiMT0mde/i+okqyXus6/7uHxUN0pT
bYQ3DRyCpX+A+Z3tNTeF12OVPp7+FK6biYg1hj+rk6B84+LX9vSsk/8c/jaKHGN1Qj58YfjXGz8Q
f0HTCl0V57rjuniQJCvKltLv5i+Dmk+sQhOUvuhGB3r51V/qaa3MuRcn5dwxsur3/7XziXR2tXcp
ywkP9rbanYYEs7g9X4zvS8rAcimx3VfG3fl4Fxn3J1i7tlcLJfb0cDcddYvjeFck/LX9JFTnrgPw
aOtxqE13sstekjEWfn1kmL308lVHHH9SVoMwZ2a5fXEUmVl3Js0Nt80jVMSk/KWXbIjQWc1yWlk3
VYExc1UCSdRa5GLBEE5l4zV08rHNmsM2pCo/1sncqzT1kM1okkKh8GiF859EwU5ZwII8p9tJDclv
t7m2iv08iy9qPqcnIlAM8Bicray+NmjQyRzuxK2W5CcwxULdTC6zkZaDOqdtChRoz2miAg8+NZPa
bOVgR0IqV64d2xFVmoK51OKVmsyTwgh0TiNgWZLNSxp/v1wbQu4KMfc+mnF99gHiyShzvesO8uPU
xtgfsfsSOMD7NmNiYFDGxwA4/jPo/EYnaacFEEsht7JcR46pJWn+OTORRVUCM4j83qWg/AixKyeo
0fZOuBI0og/bwJXjijZwtMQsSbmmKUzoeOazPcUmcO/HyFCrKLwMwJjrOU6ECFw9+S47rwDVW3W7
bC3GSMYOiXJlHj0cgww/P/+TTuRdLx+CaxU+GRMOd4lj7LfL/sEZFpNQhgAmHuCol8lhXt2Y8qk9
2Yx51MsqQ0lVBj/3uSpwsmNoE4NqJxnS154cCI+G7Ffk91JBuXxS+7c43Dz+Ticcj8glz+7IiLME
jB0cSqIZwW8Wb2MAeKhTqsIr4x8eRFpKKnqzCWt/FMOqWVrGSzrpqsSNYBjTCwPNUnaZgWWmiB+/
Yq4u6nLy0nXSU4wc1ONqZq2Qo+Bx1EM6bHj+NmmPxW9nDVI7gHZIEEJS4pkAlzt0+yezT6ujyhmw
snz1cXWDDVyV2VAWXAqgzsEu/eR5bPwoRJ56WIhYlF8GpoFk5G7h063NKFKvPeddVWefXhJ8ARzk
FsELV/Q03KrdqjfeujEjVqgG6XFS32F3JU5+p+aeJ7J/oZWQPV+m5ubsQXsVCI6P0CjY5nUKqeLa
v0HU28oJMtg3RQ5e2wiFoQulnGEWB1dhNT+EbxMvfc+3xYk0eooyWCcsiC6g4TIcH2Wkna+l4JX1
K91ABfI3mT2yB42ny/OxvyL/RblZqnWfVqjjKMBM0ChMvrEBn2mnKp62ou7Zz8MwQEcsnpfVsEo/
Hogan+5HtOAcivuAemgc5Ihxyz23uE62YpwMbkjbp3ZCQC2zUrv34KmKHsAQTbioVrEZlGO5BhYe
GnFeRVkgR/GW6GRtrAmiJsL1a9fw9AEoVeL9EKF7jCJLQGoDAsedZgmg95IhvDlfqlAXVhxySHZi
89U9TzKzGTB/YEaCZjwjeO8yajF6E8YB+nbAsoJEVXGGx3hPvc2VvEhIBidD7kNVE/H7smVoiBJE
jIto10OjVyBenOO+71NhpL5NsboI4symlpTQZARDFOHyCR0rl4oiJhQNJfssNqJDBRNQNAo4KbrQ
YNMhQ257bWEbuelHL3H7BVFqhuaEZKQq+6UkPkuNQabw7HmwzORUgH3hfOfclpiPI7TGIkg5z4LS
3yjO9kZqlNX3kC5/NKPysH/1KmmDzcAcjrqTWcalNNsGHme9AFsdInTKgEU7c+ZQ8uaAdRbjisAe
SEyfwVmcDmH7MZFIGthAnMvl0mqb9Znrz9D/89G2CQqirZX62nhTy0C9eCAVH1jrwD+Y1vQMK9Ze
zVmHnLiuYXnql/7WPbNkJY6GdN6+fEy1cLeETOCNX/HdgxhGrdUPoPNyni900sTKln0RXchdMcs+
GIlSuq3KghKyQXd4yxfiQwmV2jS69kpX+32R8g70sX76BH1I8b54vN6nwiltPbAM6XKNoc5L0dZb
BcXLcJ9aS8ah4Ppkfh3oh9Do0LqA7J0Om+YbzVIdGW9TUuMcoD327fq74P6h9ppQXYjLLRiklrY3
D/4lIIiOf4bC0I2DpxzJPjlufD7Ss8A+4sSwLziIa4hEtzC1bGmJXQsbIwx+EWu8q6To9x2/wKiX
f1s01DyYeLgEojb5gc5eOWJiM0Tuftra5i44b0AHPUHPVY3RxU6J4qsM5NzjFTeMdOp4ZnAa2bpi
3mMS1QqXRyTev1Us3J1EZtwN/TWjRG1FZaWvgKp4JU7jPaXJaCeWYelTMQw/M95C88ZhineLUoHa
QAKZOfbw16V9uvoZa1vCrgc9ITiAdxmleaUxXZk4/hztKCuQNZ+8IJwB3rT4TQWgzGQK5ldcuaIb
wsaFWUYPzQxvfLxohbAyaPj8nE3sskFdAICUS8bQ/Z2qytg4wDMVIUupYhs2bnCONDsRjKe3Zd6k
Rl5jmCqPMiXKclumMLgtiM93h3o2hpfWrGY96EwXTDdsIyQ98CzJiq4UgyJl3b7kyktrMY5Ahp+N
jNI/+2toZTzW9JzWu46G43MccUtCHGBxA6AeSPbRs+eIQy7H+JGkrp1zlxtdCbFIPNtamrprkos6
ZxyJQWDk6UKjgVDy/x7u4RAtwmM4h2TtYeRRr09D4iCBL928WgKYM9DPTIuyBx7OyOWBmH1K8Dvb
XhZYiH2dAlqWKW9c1ACy2veM9EuSvCOn2zOQXSREcGZjehmFssA3Bc8rVWhBQwodvY4bgdkxvmdh
5CjJaYQskEBeCk3JrrFXWGbGrPh8NXefHCfUROT0y89s2BTMUyEK8XnyXQxRO5Bb3an24AtQqvuz
H8uBEFD75dhOjZukKFkIzOaAKwvnrRUwcysHOwbVPZvQ9HwctmFpS4u396smScDhSnh+vSwes/aS
AmWSS0qzuh6qX73MeXYxU05meZOAe4esrr/UBMjD6H2Rp9XC6Gm3Vu+wRsHwo2h41LlteV5TD/md
8rAV9EcadoI8O5kNlgEUKJLjM5q2iESAmes3lijHtOdQ8VSe7XnEMNPxekZUeH1kebTs5Ht7aI4M
7ibK9EG5aYONG7QlFUKtgq2c0XM2iuNPmMFRBsLUx1eB7vND1X7gfnYvPmF6khNZf1j8Jvn0HPQo
17iZDtNktLJ2GtaIU07oCq2SAeCHpW6IneF4+w54qRkxm5bquYs410K6TRSq5rq95CLVxgbapu65
h1NgXzJdvBLOXnYn6ttEbKzhgB3cRsj2Bl6O2DcbLgCZbSLKZzoTxAMkihKo0r9sk6KfDUP8gxie
xY6sVAUEWEjjDmPXzrQnt7TY+acgDmelkX5LKodnRlK0gbyvH6I6oDu0sZS7gL1OGmWdnTAtCwD/
Fsvuasja9axyn+ZhY6vSpE923bztJmLM6ePgD31wIMNBJpQFkoO7R3iatOhh5geUUNvhfQrvl6f4
qrbty79VPpaAjbQxlkmGwYqEqp+TfGawUrafPC/b/kiXUfn5dfxMsmYHBTZcLm/rniHu6lltKnfd
EnSnMQgXHOrySeek5lscP5xYrftDc1l6u72yJX2Zk4LMpZUpSDTwrmSvJN4mbBRfpct+p2e9tV73
nhoqIDuqoQllrNcqw8jqjfKZo8DUCXC3VmDNICl/5V5/e2GE/K+Ye06fKlYrVIZ8ztC8OCmjoOCT
yj/rrwATK0wGQfYcJWe3ru6VQ85M0pPkGchymbW6CM42k/yKvmq2zTBzbiJMqVqza/XnJBp2nHH6
BY7e8L+qO6WVF1/7Rg2mWME+xV4bcHHsogUoCve3G0y8P+itHz7vrnNa1UhvHtowD4hlIW6xxVqK
PVzl2vU3IrsJmsqHKpagCbx1W2gn4w53MSBh8JdVOZykqd3SCGcBEN7Jx2zTkjtEV260SLlJ/p2z
LFYYSmpnf0TZExsBm9vdZDD2g0EO8o6+75mi4NFKm35kYKlOHS96hZVRAUByQ9y9cjSH/N8RDSBY
LPBY0p8XgEbRKy2nvxXhRb4C8MdgFhl++PRynG6ma/6QeSnsdAZDDbG0Q27t9AJLkoX1SlmB4Aa1
4vnCovSY8xMBa2wUQmEtd1+U52bi3JKda6IZ6+ehy998TDBj2D1Zb43Ku51UGzLyJpzs9rVrr+HM
gADzD8JI+RbzU/HIdrvelbH3i3HsThp/EEEoVI8IX+tUrexW+dX/gbkeAZv+bL9Z8OGCxzBOv7bA
e+dKsa17FcYuNsWNv+sJVF/URl214KQ0UoYFR01cgnxn3AxolH3vkK+zqhRd7lkoAkDXw5yyXKG6
rC//RRdtHan4c7HH28ohG4aWDznftvf+5KfQVF6d6lrhp1R4e/4xJg5iZjH3cyJkIwKpYuDQV2BI
pwJoTqoH8DbkHVxRBx3lwfbuMiiWCo0+3EHfpQtBI2pUWtjjkA1o+x/wK0oxFPd+FUC5j5/hmw6s
e0rTqAgGIqv1bgja3S4isk4NiR2Gn1kpmE3rQ/mzoIw54XvSTfhwmRTGWgrAPoU00YaG9DfXjHbq
XYpjuGyc7h3hGZhJkVBu8qvbdMZtXfaNwyFgxGeDT3WnP5s7w/vopb5ro/O5QadEkQmDaVTNNOMK
neXa+xSm7VdNRATLEMbGhxLnmpLRiMr5++4KPOpB989ZAIwRVDzUunKmGhkT0Yo9VoaEv3zbYGxl
noUXETkIhfWVh7+uEGGc5YXBmEHD+6AS7L5+t32lzhrSlFwaJIauYIXVkkqWovLSJwKWIOfdXgHU
6UJ1IP7IOCXLF7J95y7Cq9y72Xd2+CMTOiXYvXR0DkqELC/nzq+EVn5Axs0oRIXqrmxzumQUxxZm
9w8ZPLLLigPb06I8j4X1Uiawyfsa/ashaONyBvxG9TsI/mHTWAAOSwJsUH2vtfdASN0/4FfXG9HV
qE0ozRevt+sll8HuVRcxRqU/OeRliHnjcj/5J0EnRW6AYei5HtZWFtiBIKDbxLROEbfmbKzn+eN8
3PwK1MAlfMnsTJF64henFDq7g7KvSuPe+M/GbQDc1TG44xz1k40wmP7zxYgpfqrYbCJYm6JAqQnu
D80jA/iJGqP7B0sIDaSPfEZ+5sMYWoyQXzahbkcH82IgWdlyyOv5/qBehdSasKH+K6mCE2IM2iRo
yAgsfAcZ4ttohS8NiH0I+cdfDTI55fydWgrk4fvFt7TklkiQ0vE4S1f2u1qynTeT8/spGi8t3cQb
ZibBB6XvmVB0KYn+rWPJhIizY3mpoCoAVz+eo70XuS77jnvUIwcu+LKusTl3C7SkDYwuUeeHkwoW
KyuCcrYtw/dIIimjc6yUoEgh9gTs38BtShhwLqvGjHrATUXk/5hypVuBy94mff6h3ptczRMYVNLh
GSKGoSsGOowRVZkXs3FRmsA05AprNq+upmk5+///yFDkeejpVy5/iLpcyJgkqK1TSWoxpZjjT7Ck
Kv3ixiNHeWWBgoIuhU5XyCeKkNU0fm8pAJfDcrbQrCJamvGUJPu6uhf5Zyu06YfcOe5iBzQWwoXn
QEfvpWVlqSKkIsBwGFgyv+hEiKnXsTVCsVMv9g1llUzKc5RMbk7B7fA+LdOhEd/KY6n2Qa3sjSru
TqdBgWPcTKGfs0/HrUNKy1CFaQH4PBfuct+YSXvgn4cFdYj7sso5CkCHcQbjWp5xhosjtZghVpo7
GCyF5rP8bNaq1IjYj7HcHBpT+MN3fdz5ZrMygs/Rlvi07swl1PvyOa283w4BWa/RFkKUGWkGtc6F
zySF5eMqxO7B5VRsgRT9ANLkWwed5dV+UStgsKFRaS+mdzTmw7zgMjNiz4kaCMzZmLngbRGQXAjU
v0gSuNKSPPfjOCjMdKLLMVr305oOkYzoP05AfimV6eO1vVz0WBK8+3q03i2uH4eO8xiAFrkPdL5r
fAHnNTuTzTN+/UPuYNpmt7N/jgtxJjZATlpjfpK5WHD8OfMb3apupxJCxgtEtfHyfP09cnbWEcYZ
aaWSCNOUfW+TPEfC+esUiKf5Ko/P6lRQQGb/3pJC3E8wYyQA+10/L7pt6ZMvhMGumaveD3nOrUY6
OYsv/U/Uel6RYtkzZeQKUOuX5OI8NhUfju7TRPH6BtEUvjUrZUgOnGCZING5Muen7PHa8K11o91X
oGRnmldfMwoIbwQNzlY/X7pDGJV1SZay4iyZjcAGjIkFqZ4zaXJJ/e0nRi4fp0qPK7VmYg7tcIrs
WjiloS4KCM+ancxJaPuxRZDjQbY5opBa8UCgQpGH+3rKSTc7GHxGVZzm/QB6X6YM/Pnmto7CICq0
vZzTIS4Uuhf7Krz+PiNURpOIeihLF3KB+JjMcusKyMLinwQ+chP742+nKpaWKXp2gB2Y2OGSyYF/
z+kty9qPsKIUIwvJyQdn3SDGz6XyUOxc6WrBQggkHue2njeYDDUGCqwZoYbXJka7FgCyWHw0eGwu
RQQcOnguQlevUy7mmIApHnusEdumq1ZzVURGBY3wchziUUQnTDhzjQR8HO9C//l8+bHVjpkeosCF
LGHoM90hOH2u9BJmbGPONOHPt6M+NIasu3eH4I8tImg0EzvZ09RPiSQecDpvdVLIpHHYDEKUvrrE
mc1KHGE6/xlmoBolEJQsFYac5ye3PLH2DieJRjgfHfKhsy+YtXWypnQovt8LdocaNi/+re4d93Re
lA2skvrM9TQCNXbxgG4YqZbwG9IBFj1bOo4im7twm6G6JmjjcrLAwFHqipHZ8xSq4zi2Rnqx9RGv
pW8ja5dUKS8G2Ig2Eu6jpCxYCThEX4Pic+gb/GyDNmWSVlTzThfdFB/L43V/ErVlxcoxZu/vzJPu
PkEYY/pWV/wDgSYC7PYdo6GLeovm6zVfPjT2PKZ5CqzjWBde1VvPB0+RPFr7mlxdYZB9TiKDfgxg
AaNrLuanbn9eTn9MiFkhqEbq6WmSiwbaGb2O+dFUiUecxrwLAsleRSJ1xeMtupPPaIU9syM+WxcY
iSeGzN7JGYu2V4sPRBNnEkumVOPp3GQa2liMoOGlsI/iZk2YhhGKnf6diwXh3prjV/iUySnDiP4l
c0nHUCusXJijy54i35FYht1tb8qQ1/b5ll8EyXvPSNGijPm5dmbgdZedWKzZL/EwR+HpfZyeJdAy
+t9eOAnoxXmjapJ7Pa/7lAvBFiCiLJd6+muzSHcozeTdUrm0tAtvrRIxZEdHztxK17A2oO5xNcOd
i2xAWntnHREC7Pah6TczlwZOREpg3GVNwRqnfTQNc18pYAgWeVeymFwDWwtpscDyoXIWwDMtFmmE
Q73uAb5NF/IjQssDB8HxoPS8b2xE4IPQWZMT6X3L+ZxUHdL6Stjr2Ogn0gOlcNfMCgjrla7uw0z3
rzNZOmdAgqhvB6/+/0g6DT0S4yyNAhBnACBceMQwfui4k4jPpo5WETyUjE1jlLVV7ckWiFa4SkN1
ahNh49VLD5vXmEq6tmOQWeKDeycBuiF2HMRgeWwEha4SB4ebjE8jIaVrm8uRvbGqtZZM5pGaP/5l
S+3eErXc2QZzMbqC+o2rZsyqut30LQ41GAQtuJGlDuYHL/3SJQO4qwS++DHMw3RU9GEciCkrHp+g
Hi6Mty7+K+jcwGlAMepWab5zG7LTfqnkVTakXxGTMQBkRonxi8G/jvt1Q24k3Rg031VvoPb5y/nk
jNFu/hnOXBYXVpKD7esXVpdRSRLx+laFg/aLfAgZV3RhJEPdgrrvb1v2bXpJPSJAwtiptFg5n6nk
8pjQvwt7Aj6jSqqTYei31jPI/G9wpvFIlpTb3HacAeC+w4yK+XNEmKNR5mG/D8/SviR7CUs0sGiz
X43xbpUt34ujYxXEWhYR/axiqWgsWCper6pchUhP5ILPGPG6md4yvnxZ6y+7joK2LmuUtZTiLTNp
/bVk7u1JgIkbH+By0vY8Rfq++uIVyxMW3N6IVythRCfEg1uuNyq06rxEMczyXPX0UzEucgMPv7AZ
JFnnn9WkTPqKVFKfmaRsTyy28IyeMpnk2oVF1FkBwiu6JyR3b9fGH4Pb99i7NuFTKPW8Z62yURa/
rQejJTEHMfw9FLMdg510203/Fp6pr3ffsjELZz3AlS2qFfnYVS2+3KrcEtq6LvvZNukl1M28oW2J
iEN4USdw0Xt2GYuTK6yczYJ+G8xNn5zSZ/+AbAegZ5HxERhJk4oxYbZw3HMO0qIRXeSHCa3TdQeW
CfCL3Yl/2zglqzehENKSLnRzAyih3iDCL2QrrY6JPnmRGn+90CWWkgHPid0iFsns+AxI8r4QAlZE
poLQcYVtbGPMvbApaQ7W0XGS7FDeiN/VFI0Hqr8rklfeOXgemQjVraK4f9RMIYTn1HKDYychA8rs
Y58GRMfKcl5xgnHGhFjcByYkyRcksVNRzqvP1erFpBjwMApspy76p5GfZ5zM5N69djfXl1F/a7o8
zSYZurMD8+UiMMvYDErfF31PbM/s0uHbwSY99239IlV5L/nMZ1kjyFryh7zpf8p/GGiDqUh6TJto
Hgqig6KffN8nKtUF8Wqcv/PeG5Xpn+x7C9EBw6fjVwHa0RELtMLLhdIMeuAdKdQ0LPpJakikka1o
4umF7sFV7WKZi2hXoGlB3Q9UKIN4qZGtjo6hmdYrpA9h4ToKnWnmhchpBbUvEQdHaxvur3OiVqE9
8NIMwwPp2mUgUzC2Sm7k9KWignZnqVODmMd/7BIZf4Rt9PYntVyrPQLxmIjlSqSRhYtzXcAwdzhY
pBhAS0NCWyp8MdFLms7Gi23BfhnxL6H4EAJfKJCAjp5oTFpIkH9ynQN43qFctl0Igesty4Tj/vL9
HxROY3Xz4P+ZPRRXuOT9RoikfTqcxrPHQgIPcS3+Gt0j3Nji9axVOSqBkJrn1zvscSjJFgPrLzBG
j4YM/JVZQcFPhTZikxHh3fjR/ms4wXHdcnDG3Mm8yKxA72dEeIqhyuJ50O3XOJoeB23jz/KjEjib
1y8E+xChQExJt1CpKF+SiNmrRIoQWWu6oo0de14KPuMh9ZLQzqzvgBhcHmRquCKSPfczmVLMmrvt
Qi4H7+n3RvdDoDyl3Cv68JUjRJpTzIqMBjMzvAg56+liEAzru/+Yl4Hqa9Vvr8LluOoyVZ6DYmDY
e4NfKzCL8ClHFO5Chm/U+6YF5q1/3n0F+LDJ4AHSJAGmMK+6Br31S70XBJp9EVUt5QWuO/ti8K27
01gSqe04YdiEheT5h4BlKVixNyauSrBppUM28C6L1u1dLdx5Hqj6m9BiFW1EwRlZwIjMZbbhu2nO
8m+0pzTvYIgX42X9Pq+1Mq0LxzY7YPLtOfjmd5j1pRBnnvuGcqNbKLbXnSSqDLFP/go9Rk2Yya8Z
LXRrt7RwMBUgmw6b3GQM0rZcLIe9YV5DN/L2780Wk4m2p4mtesIPuXk5v0zdmH8WVfo42D5DIilt
CB6U5VtXRk+RIOhA0XZubA149NqltKDY39fNezeaDuSKxd6aabdjyHGQ3AVAFEOUDjE1q3hnwN2R
Fty/CuJJ5QoV8iQ4I+qcFfnbO8QkQHt3e+8x6TsjLsBzEYJlpNf44kj2WvYCen9q74M77m+wnr3H
NLi0LWu3jRyq+cQnTOPXgBVwy65j3l95X6a3hPKPR+vQrHLlsbBwYRDEFHbD8ZsYKx4gVdYpVvz8
yK6o7ZT4JhIz0Y0gNQ/3a8iYVrl9oSx9K28IPl1HKMr13Ohgo8Byz41AMWdqtRz+0RUtnMqUqz7A
vpl9f/x6kesHpozdB7+paElVdE+i8OR71ApR3T044b1YktX4Y6y+iI28tOOmOIeH+Q/ZPSZTJ78H
lqJFMVCOcsACXxetqsFztuphoAdrFc+CUzlwwP31zFmUf7GjvYFIuzJ6plqiDUdsQHWQV4bs7c+Q
3txDxTA7f/kgOIfoCFoXjNA8vfg54AAfSrwl5jmkO0NW42O3YNeItKkN+7AGBlfAorCjocjDiuJP
SiiWtrRAY6RF0QYUJs644Dsb6hDQGeT7wcbakaQFJdSz2shjaoTREtuIEQOVL9XMMZBxN3Tpnt/Q
ejslRtJhXxHcgMgR3lN0hiYNp48Fz9r1beliOTzAuoKzefWbOi3zaFxfrPvB9NfdYToC8kuDlzdS
SnlXvAz8bdiTgQs42QkhdAKJFVTjx/PFNPELStCIB0xBXP8vePUkmt25PGX8IBTmmzqNpJ92/bVo
+YUeC57NQZLBzMKTADBmphjBlc4TXp9zIMTl4+bgGUKJFtrffs2WisKvc5rR56RGfEqszRwJCM7k
T35zbArST7sEb3RGUUh1nVqQ7vS7Sll5/qZXcoYuwgnkzz5m6Cl0/Z+Qnkx485hZXpS25snxKO+d
ITkW89tqR0R7pw5Te/an9JpqT8K2f3RikhwtR5LUlzVeYy1l0RwjBAB+1gtKO6k/IWhGQ4ttEJwm
D1OUNndoqmSlMyYMeiNUUsrs678uJv2HdjQX2DZM0/FJ0Fv+cJiuTaLO1RQUzyOWCNKqDNoed9hP
G9iqrov/9r25kVav6wKZwwB5BKY0ZVGuiXy4fwVyePPgkD3SmGVrKnnKNqFsWvROR6m0cuqcwzIh
lQxG9O9cTr2mKo0RwWqXtZBwBTvod/a1ATZ75H2bVQMzzXPVQ9Sy+D3mOytU44Jf4o6VNtPODfq/
oLd+lc9g5HnzgaihCTJdb5PMbFTX0YyYXbz43Q+aJnVMaY0QhZgl15avXx7+t1bNNmsEKJSjPNSo
CQpVHOZBDGJMd2xDryDM1V4ZlBmncpKRCUDTFKza+6ElQoGVrz7VxTqVYLwZjzr+rblrQ9sb/jok
QHfcA8JYRQB8nAFl/dU5ej4DzFaS9GbFwkjEBxqKGOPnGm5Pp+gw5kzm8Ff9LlzMH8/UMN5ST4u6
RzxYZMuM77LB6z8VKJ0/cEvBzCFHJKuSBOHOaB5LR4UycHcc/p0I/X4/AqGzmmSkGeQ4LUVNez7A
FVVMj765Pb0WNXjxR9k36ZXEBSDW7/bHMGi+OGCE1atN6pZKaD7SJyKPuR71mL21Ek4+YAf9CdTq
NbsM9Bqabue5R3EhnC0YKUn+74boDv5e1FLIgn5Z6QLnQeUQzIRqMBD2OWRrUS2zl9ziX5YDRxmU
HZE2+ZEQTBc+PNQG4icbfhnI47JQ5Gx+nM1gozP2eKnNRRA/n4fxO6qFWLFaYj5r5SbxRc7rgssC
UsTDrcP+uUyqZityr3Gy3HgqNoZHQwBeJaUzOZ1rJOS4GAnUMmB3/BBJ5P5GUrx5jx7gnveXlxzi
EJz28jAyhn6kuVDID5a02LiQijrq8OshcP+nlrgwzjSUjJMJacSa3zt8R6dJ20TKZU2hMash7/Ku
wvL8W0xmlkSKsBHKOItpM5qCsmjpBB8Fqcnanaxg9v5UueoJ5vJVNrMf9VE4r5+Yyv1m3j7Iob1r
cQ37A20mA87NbkyVkpyM0Z3+AYmEY3KfEKnJzLd1cVmz4FEons7isz0Uq7r+kGFZy0mNMTpAPACf
VX4ngYOjkqTUOpvZKUbcQ0WlCZTlh8QtVdJXiREYhzocMuGsau8U6jpO9wBL3fdHpVsFRmydzMY/
IpA9yzwzECjlkHffYjeAaiJjSWQIwYoGfgyY+WUQ3jet9mvuiyXtTWtG6Xwhr6AGqymW41ipmmWi
OByA0gtAFM21RV1uz+WRGsifghi2WIwtj18/QaBIbvpCy9L9cW7MPe7XI03gbSampOm3fAHwaJI5
b3XdT0RV5evm3kyjfqYULNwp68da7yKskWbUqE06x0YIGO6dpNfxQ5UeubrS0J/Z7ec7i8xIpiA+
ToujfXlerPWWSm/qGsvjm32VDlqRxleRfn+ZVxD6j5twdl9VES5J9pmNMGugifOGQamdXEGwK8VU
2X44jKXdL6V8Mv9Xy52br11WZZD7BISQgWE6THgrwi1Zn9As+h7ETVl4ITgArkarILv8pq15mupt
2w/111bVywQcNhVZoGJhNDcXzQVPj2pzUI7eJdbRfZqU+2xmimYwrjscbR/D2MhMuXmjDLVg5mPb
ljIRmhq5InbZg+ATHC7PemN4elFiB/Qx5bupAYWPQ63Hb/oK1W1QaOzExMqzB5jNM/q56MX+jg/D
CKeiY//eOaM6ULDRKBVEUXDXVFGzcbiVQZG3nsFoHdG12kryIDa87FvWsclu5DuWLjQQC7/eJlpd
zv2wtBTWV5abaejoTGjqo9ZFQxE8Idl5x8bFzDOR0rKo1q3yrCHiYpanAGyFn6NYQE1y1JTX20/S
oOjRkAFjnARsp0yGEIhjAy3fnowPUAAMJRpGzj9yb1CWhiH/XafuzeoQJ8CtBdTUqwyIqcdLDz4q
xxVGjT7pTpkUKZSBVt4Xsn9SpfCY4TlWsg6LQUzPdG+LQEvitgOjI4sk7M2bNNLjMRgjy2lNwGx/
VEHrVfiuYLFJvIkZG3Xu/ZoBwAoaxZL+vDGXDdzHx3iySGojxauElxfK0wHKH6QAR5hfHwBFi6Bi
rPG6r4119q1ewIvWkhd+kzZh+nQsYI/kfokGGBtA9Ha1yimDcmB7Oy0R2FXqwd9UYlk3qRE3lJR7
cetXVxoQBNZzu1yzoeq3QyJY5Dw4JDhsLbsAjz/9g8WDDosquLGonlFId7yjeGSSwG2JY+OA51Oq
v9CIi/oT/r02ndfcpOiN92qErn6AgBJhz9P7VIpfS86Ob5lUwRVTqu6aFy4MH/PJTyTsjLY2vkqh
GvxbfdIIwoyr84ame+ds+3VEQJty2huYfOaDEsl3m+M7i9jEqtfGMBoayPdDTxAC+4hDoawBnwRc
PySMNkxD9kSidUXNoE8n+6DLAE8iOZRSws0stVQW28+QGBhSHIbCYQMjXWbl4GxfHS+JEmSrXm/7
qgxIAXYYxmSOT1buJgChqE6MRAhpkjkRyOYqxTaQsj7A2ekfc5oN6D66XXJkhWWRBZc5jxhpyjmo
BZ9RjNp/U/d8AtFk6Q9gfxXZJHUReBmRFAiLuDZ5rMPOYbP1nfdvt7T9hICbZXWjfCWsVmStrXV5
Xgl4W2No1laGIGU4/9BNoN/XaQKIPsNVI1YRLS5cwLAXo76xSc0+08uj3QzP/CCDwp4PrGa9x6OY
Wg68n2vOiqfSDLPLZ67zofKIaeokSaaSfVxwrMGIfK3Qt4kt/Zd0Ez332TbWN6kbD8L1NVJcby3V
yPN4mD48kqF10wMZABzIEL+gZAXdUjn9BDEnWos3rAWMGXAFSiXmIG+kfFWMEa5iwYOA2p/d5Q6e
0mjbNmPOofUgdjZIkN5an40vq4oURhgpo/tDuc/ScmA3bOjwsZiGlZ7coBBvUJPvby2lRwoDV4Nb
n5nuoQ+omFGbydBjpdTw8/Il25SwspDEEfWKSWOM93qBGMKae895A0qh0ruDjgEONAQt7HdRqWO9
1k6oTgqfy6iCWmZnWW/QjmHtKO3MHz6IXBQBQmEgpEaeHXLw64+3xXm7VF87BIaaCU4mQJBOAuU4
bUHh/eQtSzB8WIVKPRgzBoNUhEy21/e5lMFC9LnwTxdivxuZyc9nuSm3pOzyQd5Yo6s8QP+bdW83
klvonp8C1xXvLaOzNct/Kq4YkmAQOQw6DSnnYwAesxnpr4uHlCa9gnjmLMKt659hyB0Gz13HKPmL
E2IruxjHYSftLNu3oT4GOe3TOCdsDOPl5JlQh/E5C+y43oi/nlGTsFQ6iDjIyRrsWHRy7ld6c7iJ
Pslehop5FuQgCKi5eOljCof7lnTjJJppxBkNlAJJC9Pqfcqs6i6ISSzj2aBRp3bP/1nLuJqw21+Y
eePGFVJuKnSgFBCFVq1uv5R5SMis94hUZa+e8KqVf7RokJi8w0JUFGfNKU7Ut+QLwstfPyrtPLrr
6bvfvXDJ8p/mwMlMLr77EaD+X3GPYzGaT/rWiFMjKOoB+yBVLvmVnKOINTfAJsbLTuCx2re0thSJ
++PMhFT/KzoOALNCl7rWSe2ukn8tGM4g8kTT+gKWmPMZ4ZX9O5RQ7QmLUAFPQ+7Iu6Nh8BjqlNE4
CzOmqt1UahOJFgo3YqckdQmDP368jnQmD2H555zd5iMg3IfNzsxTdxXrXMNyedB+iHRi24RdjgqF
+ua/imQ2RfNS06WeyrB00jL2C1XrDh029upRlgRSqFYJtfP30gcKuzWIt3J63CEYs5eO74V+5xRX
tyg4uWq//cNma0UaJj6lHv8U9ktlwPgYK7PqARqGwsHMyBAodffkmOW6PQJqIG4jt5MYIumFUNjU
b7DLfz35yiYy1YbhXFzrr8eKuFl6XJFhDknRI8z10Odtvo4sHPtzluh39WGpUXy+mpVhAQdrzHiG
DOV15cmiucadUfJthfG9aF3NWZkrY2W3ehsy2x15k2K9EtG60pLl2jmWzbnaWGrhA+jtRj4lVKa/
WGHLMOPa6HB3rQwerV8ccmu/kXgX7bk+9zlECRgZ/6Awudc011N8zj3xC8enBz1gFGsfZW7HURTG
63QynoxTYbBCRJ+yqcCyE+son3P0/WE7sCVVjm41lnR/EY9bdy3SMIk3O/RxF/iY0XqMssPLWfls
gVpAVvyINj36YYgnCFQOANsYcMxgz8iVXPB3NJ8iqag4SJ+qPRiYkCFBOwAYaCjy9DbGCMd266Ll
BXkIOAI8777/DDLwjhVtHvucpx8Rt70ZXpjPaBuFNq/CMNufz7QnNR12A7D22ib+Y1mGKGdSA7uY
29QANn70Y8IXaRYwGufk448eAvCCQ0lYiWPxWHTBzGFEWBcVjLphxjvu7co+Fn6MtJdFYk9WjGg7
7wOnsXg4PTUAJKChWtIGOb9x1uj2/A2SBOvH4hBPVrxI/amPdNOBooV/SnayjRAGQmwzPRYR7KNW
XluD+mxo2thFKlfbPj7+iSDBqADhQL7t7QcOtYN8khz8VQR0AEDKU4mHfUclpwvmwfIxbcd59pe6
LSBTFShqBWCHNpxLg/WO9e4Zej7inDs3RiKt/0zqY6mIJ//Q12d0BM6/1Ef7o2ueOpUcIow80V3p
SOLCu7GH7rCmS6kjXAfbjj89xWowhytYaEa/tHhwDset44x5tCJsG4ai6wdd82poMYl3tInTIYgT
mcDGH4PJ2EMAfvCiF3uZmDBTHuS2l7q3UPsz18JWNDVS4CPTSeRrXrnH5VxSxaoBKT8c8XzLmBit
SXztXbmtSgbHT/QgfubvjKFZ+fMaVmOeVUtTe5UsR3ZAF4FhB71LXLegkj9iKvqvyABUPRkqjdyC
4LWa2GlTAGgFvNpi2KZBxBgS8GdsIE7fA3m5KF9nzK7k52tZgDdjBIozhvmAc0hlrNVrLx11c7Pw
9XqiPr1Q3z8U60PmCIC351d1NKeGog2ijESct/+LTGKgnHzXj5buMrnPh3OInxXbm4xCwPtbVF77
IeC6sPeUF8miSlTEYmE5o+PLstPEDLVEmZ/3eNpPlZq5bHsOTqzO7ZtqmK78UMNZqU6P3gv5gUtW
AZzG5+EeCV3/436j1Un8snig4mI5sNxb85f6DDvkzqbb+7GQvhRfUh7NJJLc8aP3LaWB5r/qENI3
XLPBdALKMZVwx1iV8enc0RlyloKHgkAQkCJz1kt7fecDH5BCh9RwHr8F4ScMG/F1i8QqJYKYTCVT
Z/+UbbSJZcazNFaSHLMfO2FuO/SEH8oe299+GnKuj5VTOthSGO+KJowd/235i4tI7nJXxYUzVNRq
so5kSPOtmadFYurPZWYue9PxcxFh/hF9CcBTq7w0oH7C8WhVVOb7/w9196K5YfGBaubuj14iZt0E
nfUsL+6RdZK5f2LJvJARCNMl5MycRxux0JTMYZ5Tz35+qNKHdUiDIvun411YYipbwoVtjQSWCdxX
Rxv+1COIAq/Z2QWtrBjYgZ/buDhmmyucCrSGmznUK4bNyZkf9+TzdWtFd90orHd33/xe5Wf2QkHL
3/BQ4rydwNPqSRU4Ehr7m/J5gaAXz+vEoNm12NdUQGlnMf4fa4BjrsKU7bcHx7q0VQEedrNl9bB8
R8OGqrNfr1UqTvWGe24hDixxP9rXEs3P1wqLM/Hjry0G7yqjmLLVuTlw+khST4qmuhZg59mx1DMn
n75Mv4XmeNqKNcw/wc829s+RSFP625sJ40hBAQfVwG8xueCFj1NEjpwIzfgx/3KsjBgrXoRG415Z
jqM32Fa7tKHAguMwNM2Sp7TLQg65CyuymAjUA/ma5KwyUwtAKBiU2pQenN1+F3VNOD8HZ9YDEc91
ztw+TOo1K4hU3wgW3sCjf7/fu0/i2tZkBAt2I6z6/Ipb3o0ZhDsH/Z3vrJkVEfE4rgb0bctOZicc
gGma6LDYloeN+9EqG2g5BechKKWiwuvt7JBZKPUkWb6P1OlBpVctRKcgBy6JvfZugPBV4adrmlYK
he/7xUXbEbKLlG7WPmInn/8Q1ZGxiLUKK6Xw5xa2bRNurWYiKcoYXM6WC9Gf1WHFP2jB0T9gU28r
LICbB0/Fdjp2MKW9HPjagLf39aXXGHTtdy23moIio/5Y5DZA9as5jDwCyyv9w2lM6Taj4J6Y78ag
pFJZcTNeguuO4nrk7VZ2kDOEAZ23DKxwytRGBh48+GDwFv67sasJEPZlRdS6Hy4OCVY6alq3hyEK
kWzcF0PZAfs3Y2Av/1nus5lnK9tW5ZmuGiefDiUp5AGlY1j26MHQ2Bwsi8ZJ+w23Jo8D0VUguZro
8GxHG6ntqk33ZB4cw3FwIe1Xp7Q4uTNoklyma81AbfLHzBuc00n7UnhG5vln5vNRcupikvqqzLHe
/6SIQnHIEoJEOj6GG/c4s3p17HqJLuQcn/5uFXQKuabrzRNvH5Lo73KoS6yytxvcRwM9iY4BhdJ9
Lyj/5CsTU95a3+Uv7YBvrxMrY5fzvNiqM920Ch+USfgBcrcX1MoVoCWPqSIpJkFZpiKv2AW7Tb+/
Lwq8M//R2vZ4ovW5PRMJqS+eGG9Lt0YnDKXEFqeNdGkQCWYidK9Cn6jwQz2wA+Q8oJzutTUVLLFb
jz2bt6kMYxaLkx8E5za2/nDIePPHbwB97z50JEOnCYDaq54Yp8b9XGT18rMg9A0BU+8aQq4k2D7e
xfQO0CZn2JOIThxeqkMnmwKy8yotj5qRS6HLSs1sO8mRIht3jzK0WgVkpagP7L+6bWQtfav0gCcV
RvDARHCvhCzdfsBkrcJHKX+lgwmQgiKqyJWJcHciVKin/8IthCPtKYIeYsiMfOkV4uWS7+iIBPb1
w4OUhBQ40QCmoSSIGcFwAyB5RgGMoynMQWOhuwHblCvxX2Jc4NS4ToF9om18xTK7fcoVPfekp3X0
FjUoOhzOG+DG3vrr56o+YM8apMh6JELJK8eZ1w+8a+gt5/Lw/MQitHATZr08cFVd7dVkkJRFqX6V
nnkc4uvvrzBol2krU5QYO9/LpBPQsYmw2Sy/uMZuPHtcHYhkFqsu08E2iHOrbnFgu92rbxTNs1Kl
xrSNe9rSRv4+aU8k0R1zNw1+aGZTyJc5wjBTHGsnDpFZaFsxmwCP6i56wpvLC6ImBEgKdUEE0oKx
ucEMmQygQkqyvgyMjr3AbnIdwz5rcWecIRDJ+E48TRz/b7xEjp3p3ZMBODsZGC7t0i4woBHjglnx
ughCfoFAJcmlUEySm+rWIqjGi9463E6uMmK5P3Z0e16AXRxLeje7L/KGhl8CyiIn5V1whtaEK5p4
v+E8/OkHhLgnczJxTOqyRNteA4GeF9OXFoSKJ/ilKi2uuEV+5/Pd8XfoAOz2eC/U6Fv6sPNAXdl3
b0QpbSgv3zghbjFYbhM5o/qXLQ9azIW4QpDw+j0tVTIYJYUMn3AdOSb6oqMAZawx5HrmIpeKMe0B
l6sld3AToOlFYIstdSAQC9aFyjhGlgyR4nn6iiuLuvlFn2fygFZLIMVKMeVCnylhQjb90MBwwEX/
596QCZ3eDT7hbYEsQSIAi7TEFNiJXLEZvkIMHrjtQWKff4tJi094k4+gpfbIA98wNkcPOa33ZMjS
f5p2T6CKdzySbGmTWm/h5uCjTB517orsjWNFLnUD7kx9eGMWwULSZUkq9bm4sTiQZPSoRdld25Mb
6DYIWA1SiRfHxRRvi3sgyLbCFPRRC0Ng/FBsfwgTHHap/QqsA+xDoOfBcW2B3vjxyDddB7l/GLQO
BJOg1ADiinyFPsi5sxMN3hNiZMkBpY8DZt3lihblNVVs6Qh0WKfKvDem0AtZL7B6K4NJR9p1SBur
0BXNV0axB4S9Gku3P7J7Ngh2NxPDecNb66GFSGQ3qoNYgw6vD5I8xAn6tyn+WFU9ltEvVVr27MsQ
D3KC0ebnD+qEBJpNcJGvGtD+0kJyLAe5Z8qqdLGvhGZ3ST6ex6BcWkOi6eoQwK32H02xZEQXP0xC
szjLFJXe8sRWArt+WblnO4YjEafR7GsRrwP4T0wbO4KdG/3h853wRI1sX/e5nLa+uUOSQf/gAABb
XRmX7TmRzXQVWD1gSPNejVDJHp/lPW3P2CLqLk/64NO0dn2bfttp1plq4MqBJ6lXaLJClCoU8m0c
c8Evyoc8E6fAPJhdzp6HPRNDHDVWtlSdHAQ079VhBFdCaTtFFYsyvQesYQ3lUs3OAFxwR49yzVQJ
zJCIGnfwjoGsmVjgVK4MV57jaPI0ioK/DkF/6kzW4AiSVaLw998wequmK5GTyfUXpCK17Jod2e3+
6nTDMJemDnIcoax8ohlyJEt8i9fs9obaHqXdDC2HczSuG+1Zg1QTazA+lU6NmJt++i/l5YiUMrzn
S5ETqDg4lmanyyo7hI81b7kBIxWD3eZDAwRa/QIO2jLTrDirxIkERuXQnEbui1Z86yFBPsZZ+fA0
xZ8KFUIrbtvdsmePjSA4lm+SbKF3lJ93Q+IV6XUa22NCfitgQsAQkNMvhICAT+atofDGXxq30ZwO
769L6rMXJGU0GN/5RpPcdDRHboeCISe9olnQOg4e2qjZNTtq/g+Gt4d0pQabhEepuQB7f2DMVmo7
Lx3e7L0yVDUkIOfF83+akoAjBrm6JzrOiwBLvioZl5pDs94vZ+w8gYift8tUPrVmmva5gogXIDcr
b60+AUvqnd4ETgSmpM58ZRvYceWg9j9jj+EWrnpqfCAqGpPDTVLzBGl0i7lKw+F5wtnP0jtH8g+R
azsdv4nIyZetbolnng93zY3d+ypH+o5SZpXkh7TUKb+EHNW//ByUVDryvjdlKydBc6Y9Lo26l6Ur
iEtD/hTlPSJgVv1nALSqnvAfQ8lKOUKJ+zHibLU4qsueVq0cNhmI6T7GfuxBawLq1rqRrAGMxD+t
tcI2ZjKcnNR0miMfjh77HFXwyiGTW0iHgv05P5VfcA+duGjP+SZmNt/qfjFsbEqlvIoc1R2DcGqJ
LOXQ05k8FW+58riJU+/eQ7eM+4Y9bxcfOslugVuKOW8ApjDBvjEe6YbFMlXrrOujFMgaEgbNaFBv
TdF8m9mGt/vkE6eQUgvU0gnGWV04fo1LByhu8EyqQOlWu98mCwkZ8URpxSh4z9xyWcQBlrgSTaMH
3igQ5IUDI9Tgl3PnDnYFZckB/UAMdbwZv0AIB90+mGtv5Rlsgoio3gM+NObDYkP2cB6JFVLyd5Q8
KM2/d13xT24MdNNfyGJEVv75ZGQ7yJBDeY3iJENUKl3Sdd5mo6hsD1uM5le5skw/5bbXRySuOlZq
XJYZLAsuFADMTIjFdWeNXG9E68JzgZq38gBZiRE8Ej5gXdM4XAUO1pU/pwfaEqraGqxXIyoimuVR
vahMyUQ3ZfOgxcLL+qBl5DtjrFHQgVbe9KBhKAfRgVeYXzlhu7mM9aUnjwpQ0FvyFzUvKTiR+dCb
JMuVv8UJ8kT3Fq6/P5QIYPwL8+2AlpNHZN1ngEWYIWTJx/dBl2R87mZDYWA0U/46YKpmahbYZOFk
SBR8WjfD/szqYY0U+5lwj0qX/FrQOr9Bvrqq5zD4cQGyYA08GCInukNBioy194NcgeEfze5WluJD
beDyb0cpGslMuHWCPCrAAyxVYD2OH+OCkBSO/b/qXTEB+tzTqlelkCGI1qj5RP2fWxKaqdBoVz0U
F3JJDp+/fIV7FZc6OiC1dS7qjgR0TLaABk2V+m7badnkZA+d5HibxvmGHc+zPMvD6uTGpBx6K5pW
ZDTL+ifgMDQpXi5NhP3FiyKy22HRWD7fHsgSDk/wDFh6zkVUBJ2QCcoMX+75xNo/d31YtGwVon2p
PTq30QLgoAp+pqobTH/Ac8mzJJGHdboZusAt0MiTGIX2rI3cmIKOZFqoktQEKVkPzS80dLYZmJsF
08anNfd3eHE7hsVl6krhrF9omxB8sFs4Foh+pL18kqfi/jSubMWruC3RaowO+PS4cOmStpAE4fmM
LDsaZe0y4jOfHa4pn9UBGgD60BZxjOcZMbF62Cpw7GkphkmTff7r1rlx+5K7FcLUubp25kwZM7OJ
8Eo9XpcCFDhu9+9RxpJ9RA6tIX4Oo2+/NqNe7ixNIw+hd/wBrR4Fe0d5irMsEIt2JR7ITyg3RXwl
3VYTfbIjt/UNnY7kWorVFRJBfu3x/zklJ8r+V8ShMRfulGL3W96D4Pf2K4umrYE7GMEvG2UGaWyK
KOkHdJgZgcInXyfzdWYWbnuPw3TZ7Iv6tq/icGPR1bu8vIiXDgIyCiv9qgwzpRDCxrS+GiQxDeOs
rx/JeDe/Xlscu4CVMbsdrbLPp9PFhO8bYUyflTk/CQMOKcsGKXrZt9FjwoLn7taam/bR7yj9tvP2
a3qTUc9rQm4RbTk7GKsMtn2Lm5KnxKQrAKpi2Q8esbGuwi4PpgDUd0Xes98m1NaNrIZN7r0wRjrG
piRVAK2kwZ4d/3CZKFVuqdBYePJXwOvcXTxtfv/5I1Kgbazail1o2NxCK7O1EYTS0PYObBNsV9vi
ipLQeXMR2sa7inczMy6/jAbjkJkH/FeRoX9lqnv32wfgBjBpPk0mDGcjZb9osluJrIShgixOiSzM
6mtnd4UWXchjdY1TE4OKwUF2szNcInJkIxJ4j3aTU7DBbKWUxFZ/qZD/XkuQwpxMVGUl96xfM9+N
z6RgCj4tNKpwpaulqzzMBIt98rRi4XypnbCawrFzTOlSAxrg+szN2NssoTSvNRLKRfTm4Ld3cIJK
AwGcC9AXgQXILZ4jhDX/0MEHlxoYJ6+vS6acW/88liZxKOlF0p0mZkaX6Qtbel6dQYYAcq3bKOcU
4UKe1ISu19k6nbq2sueHgFzZTCjJbViNvxY4qQVblnYr08eV/S8TH+D/gziDlNDF25L17O+3Pq3W
6PlDv+OKdaN+vqUAJsw9NwmSpd6IqD+J3ArUWLRpuRZYqomJSiqf667c9WUfCoGnr7e1VXWFa6Ji
vS2+iRfRtMGh550cKvtAri1c/VFv80B2LdFHH+gnKAhMxSzSALfmiDXkMqvhA/NmIj8IrToVmwFO
jqhFGoJi9XVyKvb7vhMUEaLQr82HiRRzdlpBwPdEp6lfFvEpvBaYUYsRJkVaXiWAKJpBnsnC+nE2
7OLBipLotyIkPlEM+3x4DBuTkepfHHTDeN3hrT6SoN5cuyQPDpt0C+DQxy9mDEFkMg7HGjAEADQb
fhynNQ32qJD/4nSyIb2R6FJInS1/ynaLJ26jsfm7FaQHtJazBe1qMPQoAIPHPxGqUh+/tqrwnyg5
kanFUC4v79j4zfKYZqfJ/Di9QwQCpB56hJfP4f7UUL9lDBeOOA1MUoTiczwLil9jGAN++rZxEWqD
tG3yOQ8R54XtKEMQwnmj8K54VRH90eHJu3NlwMVeGc4J22Si+2XbQwdfIEa5sz8c3gVtunWSlvSw
ZRlBTWLB/zap9wNP27lFLwRiqFNkMScdBG7sOOGAgisBsh+tuveOsPXTXfpDmYBZ2XNzcKIS2Wh9
b3HWVlOPYkBo6KoDsqmbQt4iVln0jjPTXHAbeChnRIUyn/ugpbErLeh79eVErXF83uev9IqoTfsH
x5+M/KeHD3H147o6zrXnVmg2jyGKsT4iI3kEI9BvPTX+QxjWriPfrGb1CJxo5zR3cSoqxm419NNv
Ttx7jj9+QdoEsGTixuPN8TXHUGoucYYf53dMat/yQSTEEbRupSwvswclmy7S8TbJTASmbcBD2yUV
yzzybZZFTw+L0C+K2qobYXfQtqRXwnFfyk7fGQxXm9iv6CK7o3RxVlhFlNAtfE8NpoemvAoa7RJu
8w5/RMe4B+tl9IOAvpTxRmzcbuVQyb8dd0c8Ios5xbJRQlKN8PhOqmRNGObjPZxsUStw+mI4nVAR
8swviY7dK+bi7glPT4k7FhRBDyXjlmkiiCrYCpUz2dK9ph+FZjpXI1SX12WXi856aWyHeES/dSPr
iCj86/gWogdfwJiMcDjkvVk4ivIZo8t2kCQet4xYcWWuC3K0+7xHF73AAxPTNAa6msdoqgVWxMzS
ReMD/RRRzekvcPJAd1n2nKzhmoQwWqtmynVHqZTjdQkkakLzaBASV/YAQ6BYX2MlAC6Idb7fIKfv
rv485c3xgvBWP6VcyhhYmpKML2+/ZJm9HTt0juHKFvTZ9hk2G5gBpBa4YfuplZViRCiQphjL7V9O
H33BQzsGYs+clDmSU51fmsn5WkM/2JXoNkCeqmvM4QFkKp0brp+i+4IYy6DDKq0p81hBNNcXTB1j
nshB3IygrRL3dXNXZ/jLItYKECOlzjcq04bx7+2EfUJ1O1xMBpulXmmmWkO6y0U8i04g/0F2EJM/
1fG3LOlOpJcfaPLCuA0WFlKI4S65+i2B76U+7p3ov+keyDwSturexDfrSihyAIfv/vCIFrRDgwP0
/kMxCizLY6JsB30KNcBJbSj+8FNRuxO0U0Los625HGIN5Pdj+pK3ghjBg4AuFzc2gx3YBvgwtgZ4
F7eV4y2LPzImAfa+fOQAXJ/xE/SF0XLv59woYZUtuJV4zeNjseyxARpajOFTG9Oax/MzLYL8/7SV
Z1XJJIvYeSXEBW7f4X7vG9WYr9U5EkfauFflZTJZUWMp3Ep0cmv6Akkug/JmXhVf+sgTd/Cdktn/
irn+IpZylPAr1tup53d9DNH6RV1SkpujNnTxi8M16TuTberysGsrs6oa5BzEt0MeECrg5ILLibOb
2hmRzNSwb1EqCK1kXzm7fy42ybCjU0mTTvh1/sRNCLqlOWhyvYhyVm/+IX/0+Bf97OODhkrEAv5W
HX//3msjzcXNO9PwBbPQscZL+bwQGdJSGkjp4mIMYdC1nzUslTsbOVx7boZs+07+R3slZeTKkZnP
GeC/yANyxCF/SuuPGRxy35wwUQ2+FUfHYN7whTSEkpyrc3vOT9lOmCyIMVGr37dR+nnGHbb38adQ
yybtKqYjSVGL2N5lvCrBgiBJasa0mUcKOKxGFDJbWF5JLIjHUBJlGYXIsSHAxLe2Y2F0jYAQs4lL
DwbKYoIjH4RGZZPjqsLO1P9vAB84pBObrnrS+6qvzRIzhtj60H2LOmRl9E5zXqs0NSJrva25/a42
xGBG9Ye5IWoHzlUnJhpURDNpMY3kCJppm32Wxcdawg8Y6RyjuZmU/5XKwVj2bfs0ushPb/KU6aMq
jbMvgljCwxpmBUZFsQg4AEb81SUl37iPz34yQYDYcYKDyxwuqAHDcK8i5r5S6a75W0PDKAnZKVDU
sTXFF9/OWNwyI17go1NVDgRbLsGudZ2FHDZny+auVW71ZkF+fAjszsRIC6w8dc8xSjaAypUDay08
QooEi/Co4mjLC7oUXawfZXYP2dhb60AUsxOTNSIuPPmP/Z8yI0Scv8J2tI8p3U32KETutlbTL9uB
+Q8IAvqjXy1daiWDgB8g4z1VIpABooGza1zl3kQprzNJQLPXblIGsQD6GOPgy9XSbOWWIyQdaOMi
mSwXJmV65olLqvi6JK6ghRU/ohIc4Z8FNPoZ59x7TADktavLY+tnfPEnn7N7peeh/wQJQZ8rCVix
KNj4TiZKcg10MgQBSf49SrHB5dXwJ+FssIIZIRb84Lee3fbC+BGhc0PsOO8K1mHlCUkMkPLRAshG
HoFVinnQewO06Z4/000FnuDI8kLJaYXQHyW6OZyMSbyYgHMHKUr7qa/5HKasZS6I+hGTm/swC0K1
hLID4AJFo2CjZ0lZVu6w0eiLR74EpJm41zWy+22mOfIgurRlHdibICCmb/PxTWIfPsY96+zqnT4g
HuNuqFS4QnjJjkSbWo1A/PVH+JfDZ40mxdtRQi1y2SmdHnbSU/P/i7uRR5+ja3ZbMuaQKZjpvDo1
BgUViSJ5bKgJ0wjazt0QRlkQGfJiGYP09Z/JN4cy8QhHvP9ps5rlJ0EEE8iTsHW09CAXPfXmd6yb
0EEo4MNfWhN1bEUakewst1c6FbcYRa9tHaiGru82OU/ANgRmQ11GE8sRWM8WG+a3L3oHxHAE9auo
0ixzBmMUt/SEpyIQksJAk2O/C8jhVLR+jRK6l1JNaQb4wjlJ8VHqOWXtHOtsMQ9OoTm1KUMM9TQx
PpL6Ovxe01yWfZOWAAyMwjNgemkT9PQk9qg9hZzuk2M7uBB5UhIoxr4LmMSGr6t568fC6bztiU/e
RCRqZGplltDuEqbj4FERb8RcJM6Ynuc0eKzN88484jllHWSt86yiSdaFXMsQ4Z0GYpNEeZx+4v0c
P+iqhgAbsZykA6FA0tNfLYy7IcxxzA4EY0LknV5hYu/0tQvumc7MPP9/ufv/SG/k7elxOuw3shub
rKxgTQrrj2fFtDfBJTLK7F/eS1/neuUhdgDWqcf1ENKnxMNFafsWfvW3JXxAHjCPAu8vgxYu5xKP
yOX328rqfPlqkS/DuTDBOrXbubiaaO96Yqz455y8upkQCxA0IyVEuR0kc1ym6uAV2ju9zfJRimFG
KIjKKtig6IHFAhEbncPuO/ql27e/puI3biSH8s/kxt4UuQ6aY/PZwEsQRM7OdxSVWfIcQ3xR+3jw
FsNQIPom5+Oq7zrqijPMT52Vy4FkoKDWH/zJ1FoFSX9kdv/tpREUMqti13ODmQmvnyIzn+qxtst7
wIStM3FRZruCDtvEDZ0gv1DIMQ2kKPqi6y2PfOPNOciAjmgE43amrayvNdlKftce7zKChpeJpudZ
W3YzMXQrSwrQbebp/XW77kswnd21x1+9/+Khl0QP4ZFu8gdTAQIlRMVhC4m1EU8xZeNSBSqmQQNK
Q+QQoyX6J/bFmoXdaxHBF6Bh35SwkFYzUxJ9kh/1ly2QOY2J31WCPZJkCth+hvYCRZl0nzhCua2d
MYitm3+IAwC6kl621Q/O7TUi65fXMPaAhd4pOxcONg3AJV6zXRRbS5qfvKxw3fqNAYdGTAXLpOGH
HSqLCPVepBe6xfB4koSjdCM4LKUOWm1EzlVgqOuBRAsh2KBRUaPhH4O4UOhJqA/T/jBpyUoFL7Pw
c0kEpKfyujQU8kLttQrbBUr8sG0ocAI7FyoQ9hwyVAjTZm5O5qr+sS3nRndjBO2cw+uWgSM5FQ40
gV8n5wNv42P92OyFDwuvX/f5xznHCBR0BnpsPyeuN/j2u6G8N3JM+ye8XkvZxM8CpBATiKDhHvHj
2Xx3DtjzqhoTnTe+RbId9FUHAedE2mgvLOQmS7AJ11/DM52nJRbvKgCaU/XolS5XTtsJ4DNuCIcX
83mOORTaBNvvDdWBiSr+x0RXdIvRNUlmpEuoRO8q4fep3IKXkWGBklZeV421VJaF1BhEJ6Qt0zXm
NpBpEcodgJsmxA8j/1393GHOFDcYUQzPme5D7Lu0rsFs0zwKNsxerFPEDq2modXvZILVvmoafrpj
DHwRzAy4Re9s5lTEh2nHcid6cdCls08n7rq99+jQCNC2KV+9PVRnrBbRWSjtutub5R08nYhfmor6
EZI1tJWHz12MOYMaTLa82sMgIHFXW1w5bEJOiLK2DO9jf1GHI8tsvkZaj+Q/jxo6dDm8zWrbi7Ts
q/iBX5UcwWJd084iQmRrBj5wBto/As9VUC8cluLt4De6vdxcQ6GptJ7MWAs7N3gfstHah27jls7I
eyCaUfpSz/iN8zOEW4K3Rl8N3ScNdJQnu+B/C0HcubAOcJkVU5xGRAGpDu+WDKts/j4iPHxJhPDt
PDA0Qujoz6pDkEIcsoEj2D+SBB/ZYDyAEmsn9vPkUq4SmvB28+AzAygnHl2jJVOJZ1344F0n3+vk
EA5kUappMTtAmAkXMagxH+sgiUy5x9W5XhGacIX36OrIGFaEtiNDJmOeo9sAo3PSsuZeVowqhnPG
i+Zive5oJTz9xwrqzr2hdvybQcKT51hWLVeSBJyTCAskLJdD/KZB6+mP77pyE6GU2oUSwtSEWlSD
s8r7YRt8VnSzTpgTUo8W7/zSGyBW+OpbIgzxebfU/FSYQhxLXKvHjybvxCPEt21J2VCtk93TTFEF
Gm1WAUMec4rEjoHcCm21+FpVOU/sTw0mU4bKZ55V89M5nKqfNagJ6dPI1Zmlboxqu1VT9+1wduPQ
P6ylq1oNdRLgzpe7qRctDp7dxkhy/dHGsS8myRKSEpNhFfA113KdUo93hUjWXf06vNccma/BoWj8
LjWAAwmIIAS08Pvhy43wn0Os/9Oa8lTLoB+gR3SNeemhBOAK7dEQ5k9aNJQ8c+MIRl5Xl2uIqQ2k
mNKdL1EMl0KqFN7gW4Ao8dNj4BuzoTZFtJihOILWtTS8KMPU0bUtsop+ryExhHMuxO/QDMkfO90E
tvC299AUjGzhjOSqZe0MNAnu0Mm8R4IRYt/rh8PMXqUAu8Q8ULbbj15llbg+myn/22sCr4giqPMQ
qFxHCQrMOThLH+sFxfvmUvWTn5Fwni9lM2oUDHS1p+b0PwMhsAlqLIPFOvcozwJJTct6QgqpVRVe
j8NidbPmuhhPxpenYv5RNpfruzZJ0A7KjOxE3pGXhWoLEJf0IkmaXWJIrzCF1XH2mMJhZTJcYjEd
+J0aX3/olsX4HZGubl151C53Tq9E8Y8M5Fs9nZGgzOWeZMMSixWnwPI9buygTNWH9RmJ4NVt2MnV
ux3jhnuu1/ijsNJQPByEw9a+8OwUaYeHYa8by/aiwZjkfVMqNe5UhciIwwrLksnP6HDK875x91Ir
P1OTmjgMs4/83XkWuPZEIXRZfyG5Fq6MUP/ClR0YoHpV05dC/9IjQDTRdsv5vSC/0WJlAAlItqbK
B4249GqpXlSB7Oib7s4TBxCf0G7go4SiNDcOq4POfuF8V7SGuD/IjVIxDHILXnXhF8ukKC2Vrqdf
vkXaiVBUCW9z172AMsy93KOFt7O++7qQPT0bkB6Qx6MBTgHYQL4r87dSzKVSBYLnhwEWjPBsMaHg
68M5gyPE2MYXTUDPrWcmDVnhhHQzmhHt7QbLde/hvb3Lff68kJ9BYObHs8hawWLGaKtRym9Txv/S
01QyJneT6fkoc4UgwWS5h4vcDoWQVM6CXk+qg1OBmVtk3pUZfrtCz0JXUMxcWneLq0qnLFluXgJB
5htuCG7FeTD5MEhpjLS2XH7QpJ8YceJbXFjy9hDIX2gIAsuPuk06d1Scd+KuchbBtUia+MPQNwVV
MJcAho/LfCmZN9fOS74nN/UxbqAzJxp9vkAnDMtspl3JFGMQ4deDo4RhK7cmALaHcXdfX8VzltJB
Go7osa0wjICLk0d7MFKcgwxVxfReqMIxu0XXngcz3wIw6iRetT7Ml/vqHuBAhDci2MVbfdhiaYgS
0LZGSB0gQTuJOzbBKr9i83WMn+jQ/NBDK2H7MYN85MR/+8ijHPzGtLsyYr/HzjE/JvHuytItZK1z
YizYX8ufX2x6oZbpot9F5Iy9MFuDQ9XFK7ySzhpJaH0VnnbHfEq+Y0NN/l+rnHSiIhN01/IjhmgW
24qimn/OaCw0scEGAdbkFz7bJ3B8qrKXeaZJrHEaqTzMzqJMjjqxM9UB8U7jxL0zEYNa35d2J9Kg
n3j2LIpaVckoSj1VvreElQOgg36PGbIDlQVhpRGrxea/4l5EwCeu2cEwYS+sS/sQfceIvMcfNPCC
MzHGtgFbB7l+TpSri6Ur8VHXEnuWfy5VEV1BUzMn00WsVbS91ZeKPoEcTMcZg7TaJtZ5joPMHsI6
IJGQxgqKooNYCNFQVROQmhtwYf41NxBKPrF4DPcwb5WSnyqoMzL18EBxRkOjs6hoObRPbpUA/Ngh
bS5pB8MhTTAtjLnE4x8GC0lW/eERLpDnNg7zzRO7A/9e4EnRU4P2AlWQJfehRoDufSaoPjUpJbca
lySu65KFddO4vUnQnE8IbiJUVqUQbwICUciZhydLsZPrLtaQU4aI1QOy/r9Qs8+f2KQ0HBmuH6Iy
0K2bfwZBB3Of9gdl5uvphIM+yzwlzm1NNFe2sX50N4oXSpyBfpaswZK+Q4RnjiXKOnJ5MUG1Yq3W
uQKzs9dDLnqjrGIHtWRVqgWpoYKXpEfgnrWYhv0DNlXJerBw76l3CZa3TZh08BwG/7glPn8ut/Yo
3tZwR/EdNxH5W+eXQXwA86tPhImh3IP4fBgqhabEIaycl3ttolPZAtRCV5/JqtzurTsAUJyfZ48J
4UkHjni8XKFh/YhkOc4/fGri5ZlvWwH3xIpVLg9+Dl6x+HoUuqBURjwjcaaIw1BmWkkBEfr2vwWd
f/bh6p6j35UFQyK+OyerPe+ori5xepx/oU5l8RS3TkMqG+nIfOG4upiGROJ6PZa9q0IYHGYzTbCD
67pu11DyWxHphv039aAcDmZZroniiUP5pDlx+iE+lixTCb7ICbGFkdxTMeh7YhOprcoQuwr+3NlJ
dAsq6MXPAX4OBJr4sb2R8Vrk9JPX7Jyji/yeIFlTc1WMdaRNVUKJvVMaZFbO7/42e/QiatMgaK5E
jeSIFClC85xGgJ81F5gCMAIfvDn+xFbQ98g1pboYOyMYE0HBjUOtl4AWbUBdxn+vx13M8u1Qk3mD
5dPDTIHLhoJhZPrntjwASQreJ4IDxKu3pCilDZYle1n0PNmuOQpmtV9j+1T+vn+8tg4hSQ4f+n4+
xU0MoQbXjYCoBiv4jTf2jnyaqPYpEKR4Hg3HryExHkXuv1ZjV1vbf59F9OJYCWxemBk1l8+PsNUu
ETmqxBvyvgtAXLcMV48YN8xbVA2hzYkHVmV01ioiA64gBnuUi+pquHEnsBZOrrNeUNkCSPecb9jE
k9rLSFH5Sz/RhwSdd8bRhXdcZnfiSODpvqN0dBzQ599/de6ASjVn5sQpht1XdUNmCoVCD6NTAE+Q
H3gRKZhhQ2O++3yp4pYd/J1mdMZZCZyNHErIS9UqjwlStYyuRGOcR3ltAc2ttySw9Gx2xlXCsFNu
sJa7GE9L5oq5ZqtBy1dsa85aSJxeq1Sr8OJTZFb5dF9kTvILtqSU0p382XpATU0z3a6Oi6BzZY3H
lTF2VvIf9U7ywcPqF2VBHqAj9Uo3N8Bb2QCbJcEurm+FW0LRGuzAo0c3DwIzzU/WRwnSpNwua/hi
V3GUSbJVXUqsJgaR81ERRuFAei/0YaMbBEzKwuiG5A7PpPTBCgNki7IYPjX3z1t7Le+cKPJ439QQ
hYK65oNluk4fZ/fWWcMPDN/MQV6rtBZdxcVXgkY6NVoWla7X7+9Izb50YaHFa1lHtcfkl+RFcr8C
m2BuMbxfufp/8i0Jc5g6kNNQlZr20O4tKGL+Qrect2bgM5lHvRvLeZ2su9XBgZiBRnZPCQcUHHvH
YVWSDZWlmqoCbkNfLu1y9HNdUVRrC4N5oa9VQ/E+C6vkhBA4BPBsZSbV8jUpdkqS7o6XrOW/lOec
+kObIIjg3fotA/oJAieDA2hs1LsSdrnhM1xkeZDKToGbhNSrdiGkRLwhxnbEeyjTDylH1AF6D4cr
eSKtdQsTZL1W5hWuOAEGUL8M/l6uQbG4isNY1k1fwaokhlO6NzEDWZl4PKaM02p7BLBVaJuVEP9K
Q3Hj3qM3VV6lPVtbMqPGFLiUyJgbTRidKwVUtWBaO5Hin9WS6KKRJm3gv1v6K+hQx3oIIX8OrXPc
2/uGGmFZ3rCeVHEitzOwkIjd30Ohhx7WHWPJia4Dgt5BVU5ftIvAHJ1DCT4tXQj7i1d8S5HKkg73
e6QUQKntFUYN6w94iLCCRRh9mRaWnz19GpXeQloqMHOqmDbM6zsfBxAuObmJTNgBmSmiPAcem5ZL
r82OtWNRM2lzLlnMNIJ37Avu1RwPWG1l1agGC9pLoXBjN0cRiWHwPEN9MH8bqjtn5xtJNMlpGiFv
Vn5/RHrA8GoXTs3NNbiC3HhVBtTOqbaewOidDkggJOEaiYc5V6DflUvP9sx+sg1v3x75xROzJlO/
bti7iqcib0JSVuvSP/RuPiLtherzZ5mF54SfW37/WcqHvjmzdS1uoOPT5eWzqibOerP+nK3ebt7K
YaY5B8Z6tHJqIXPssZD1s0gH87lZRdOeeDhyKQUtDvFooOBOdykb5dW2UJIaeoygmmuLODmZkHNT
A73G3ZKjv4JDtxz8OCK/DIaBGlQseGVLCjw2tV+uKwETfPIXsFD6quzN7Az3szUoliYZdvenmar3
NMn6/A+V8F0AyrzGSPuUcPw+oC67st0c+EdJSdMAlhEs8et590rIsPNaZw8yTUeW0P9HOQYMfjIR
+CLASy7FjyP+Eopgd2nA7SSy/KRSZ7JUa8I8CzBCOzEAG3JfWYipOcw32G1UsEYzZ9vIFS5YSy1P
pRrdjV9UaukciWgnerx+nyaHf6Xy9OiU5qGywlmNil7cYZmlo5tkTOSgUu8kWFS5USEr1/m/Xkmo
jiNWdDl3YB+zpxiunI/LonI1D9ute+JpElWVB+fUJKyyXtRQzFlKGw9szaMPJn+y3HC5HEcc59sl
IPbirj2jShBA782FJItD63iVxgPJK1MO4vnT+irGoCP5SwgABTePY6HH3nTFpyI0dDzQJa3uaLGa
e5xFLPEDqLGkybw7BSsX37HZM6JwXU0F81tKOln3G61Rye6BwRQVBm+fdt2gzr8oOxeQJeU6GS6Y
zt6MeHwNbiCoivqrNxlWoRZJZOeSw9N1oFRWw3Yq/Jf5MT4S0B5YTGAAxQtZIJvmoXIOqiCtL/0W
TGT+tz8j63gwuFqeK0T9km7Y/hkoyKKtadjp2ZB7Erao1B2cZrw9fyg3RfIay9WYNURp5nF4rsjq
y+e6m+ZLgd/apTBxQ6zkNTZkvqKKovQlUMngrKoM3SSUbnAXbQYEzndGoJCQioOH0mHtu3U3ZASb
9Hr1Ahm/I7tApwlBMU7mlfzNfSgLwAflxQzKpeVjHxoo9JVxcdUPAfmmjK36H5VNecOgOHgs81WM
NugmGzgHEnneY/bvlyDn+oi57KAlY9B6w+BjbrG0XtsolzTdMtUGgAceaisSCFow9YVnlvcMED5w
isN7uDP4+VK2WOK9BA7zGirIwVoGj5w8Vo5M7qN5MFk0j/TXSKSqgVZpPkQTJnZAq7vwPtK8kozn
R77NLehJXF9x5Ipy8XXaUvNG1ebiHE3wW4pNIpebW2alOpnLIdnYG/nXlhv5SDcAxrkh8UezYAnL
4baXjOCchwytF1WE8QetQHeAC97+Rj055WRtTpoYo9lSLlVHMhXf1NsFRY97b7NVYO5+fAFCNWww
XpjXsTO2n/uf2fJRhhviJLH+KB5alZe6H1G28JIfaEqPWVV7XXSMQFtjutCvkL4u54egjp3tItOA
CsRJwxoCStYJlWEeLRat9guOViZjMoMc7Spv/QBhtAN+Rd028LvfamSWo9k5EENEvZSU12s87edC
EI+9BV1r4tSyJU6tSwRWBtJe1hWBZ25p0nI5rlLo/bqWoRV98bTqK4VaD0OIwVD8S302k/QPFKJi
5lxsjtakSn+X++sh9PuONogvtnvCEp1OO7wHicQXVPNyREvZIYcQqSp5Pa4b8gSetJTiZNlb0bCg
rGOlsYEYi/x0U8azb7lVCs1xRO6pHae/PjGerNOztaSGlUFc5bJdL4JwGl83jVlOBcxfG20JAFL3
9yAkIdCa0CATrtPn1oyZHH0D7yrdU0OeLkMaP3K434m5NrG6QL+329/2pAjUhPyZf677VWRKwVhO
w1kB1k8a0iHAi2p6igZKtz/P9mB/SqqQMXEP/eXqBTiWdpfAvD3wMTqSqxw5OQm6SgATYwHgqd1G
tlQAZABk6YSj6YjuHjxVr8P1RcZJYZ5c98StaQlXk5Qs3ylrWmLlZqsqi55ciKJC9og/EBftpDXL
eavcIq8bvRH33V8NAG3qY3p7OTblRArJ1vXErlqNKxHyTNH4jgPrPlZa7R52JNdCrMPKyaxw3Fqf
Hp66v40+0eV/IQEUgvLymS2SauNtAcolAErGoqr3WWFeEeNhXMW22zsafkbqq9x4+BqivVwhfLVO
Vj5x10kbLLftpP/oGxUR2eGfPep+bYP1nXnzQG/yz5PX+m20SziutvXG4RB7CAL7DoTbyhBr0dyk
3tIZaLXwDQDm1EOLPYmdHtApnbSb/XdtkBO6AmLnVZ5y6e01DN0Cp9LkR7b0Y+tfP5yz/zugt+db
aoR7PGshiSWEKPXgXOtFsKdVrUipeH6KRjsqlmiXWS0FAoYGcYqS3y64dCgIhWbJAJwlRkY9e3fe
5mk88IBqLQhz35ifSQu9iwrtKpC1sp8Ev2A6CPSFWB0/E9s8XSrabjFU+6J6Q1jNgx8NAo3OUSGL
hG9Dz525egC+A3RifvqeMXyGzqo5v78l9yGVXvza8CzCFRB9GiaILmxg2qeNfOlc9XbRB8e2ZrDq
QCCsopmy2PxhVLMQaii1cR5OcniPvnrdU1oLdNticKgw93eylpd5ZT/fz9MuQN1pFOXxXaH1rb20
08Z38YuGTOPcLAOsGCUed/ezXgI2HZ6AjON+bydg+E5czfQbC7XTQrbVoFlZSPYeUXEmy5J3fZMp
xIKsEtSDcPxWIh9rUhbxchvOFWUt5NiBX3kG3npgmcXOZ88rz4ivRCZZXAz/dxe8vShP/g/K7cSR
nBKCYyOBqINCd1sdExHwpkH2aQH6J7Z6pnCDiootmsRkgYUhR5V1chLkX9I8WM4eF91D0nU0XvQx
r6rVq1LtE7UA0cZfo0hZwyM9fFD7WPPwdJgi0PHKCtiTDvcxWNNqg+kgHr/x4+HeGzrjNBiibVti
j/0wa75yIocZNmo4i7kH9reoDXPuVv/H7G+YyVYbrQu9L1ty2o2wAJbIxYSdfKCXbPLCeYmASfyr
Dhye3eqcotYpzL5h/qr0P21BFHwAQREdktNroqdoSwt2pTks3J03y2+MZeEK7AyViwkdAxLrZSBE
Qr1tYJaRF2Gdlpioy5UT8MNEFT7+BEtQ/2QBcwXLM3EdqF25GOCXDnK+RsTnzsOFhtXU8E7eRvmx
hGBwWuZ+Cghe510CiybuMh2ZsAyOY+vfKCrNShaptv3xAw6OIxZ5jHp/Mm3lKpF/PKuIevK2Xaov
cdJ7m4+QnRJRLgpEddF9xjSus+MTexzclaCF5+q1JBu/Y8zwwN9K3Pcxmh9EeYnxKOrRbEZSXlkd
RJajnzvtxNAFetCiH4O8XnxTxcJfZ8bazC0v+EV/Vxaaw6dx+19G+paED3AQDowSrbGwmS5lv8V0
PvOrWMMx388YmsGFHTuiU7LPBam6Wo6UUy5hscVnLABDpiAINIbPjDbzKJ8ZK6vooCFPgOofsqwk
GhMKFqxYxkQOiZOEVshG6hjwjfGgA7Rd5ig2U7wFWq2/mh0h+2n+NHmcroqfg06h5ct3oMKOvuPq
DLvRkLUrvPdNpAny8UvHTMOPi03cNj+6t1oTNVHXNlGZtOvkNF92rU7UNfj3X4M8p7Crf3uATK6S
8l1b+ts3bsolPx4ThqmiqyYIdbgG23iJfVxZxUo7f9aVJSNVVO6bxe3IQtLdYVglCvzdoZeqeOKk
TbVsimSxTrBlf2t8cLcNgJYT/fv1eHdG81/h5m7edwkxoUNZBsU7a1frtPdv1oJF02rg1ctaGTGi
FrGl9Ysc1XYnlrfUvZa2vJRcH7dP5jfcFGrcrRHxTv2wXtMHtXiwqX2AJiyWz3I89j94DayMxNfg
9tlVIGdBU0cgiylCqA1D/0pEKMwPSsHH/e8N0NfQSolTIJ1/yQKaccjd7DifY2e7B9EhnUe9LW1b
oliokUAQ/Lz6geU6v05VfOqlEdQnyOrmrEQ2T+tzeweWH1RiyyDf8EL9iPcneSmh4E/6UrL39+JY
G8oAOnDiTeSlOFgJRzDDT1Utn66YfnGhohvhymEf+A/XANYZ525VUDv+U0eYncunyoyFKA7OE80T
uDNtFtQ/xyskI9ym8J3fB/uPi60Kmt1ZTS8N/qxAEo5SBpuLTAXEUz03aiwL5q2/KbWJz5YRsQ8q
NShTx5qci02tdbonyq81AHOFRNKtllEJHId6jlBTho+GOZEpypRDHoQlci1I4f1Q2r7cNFm7sBim
DOcDMjqMh914GcKYfACUAFDCA8LTdmr7pqJnfAc3q9eTt5t5lRnFVUYiaVLRy4J0j2J54s9qvuVl
7lwCKl5vVQklevt+8Opj9O7YwOSJ8cfEce5dkHPsLhh9fV4hCqVcs80AVF/REHB4uIklJh2u+QNm
dmzsilCdkujHwOFHWK8FMYQu7sBxKx88laPBAWZYeWn4DJ4xeiaL5RtueXsW/L467sJAy13VeXjQ
aPxHWgTYYGHfYw77CZ/AyIktvzAUxGuxnS8SENFjQV2hqCOhB9VStD9FQSRaBQLTt9GyHJjV8fT0
e/tIi6x1DoRvTF39fOJ91PSqvTefvFZXAMaGsMkcY6Vwkl4+WhsKxEmK8DuyK3TFZt9Lu4MyiVhc
qz6LLyy4XahqOWvPbMabdHyxiXN9sO71L4Wo5LmeBMdOc5EvlrjilZPnHldrLZ8m5rjntDFoLsHn
nq+1Kx8R9BMWTVC4XEOgo+N13iakToirgw8exIFMxFNX1dQ9sOAvGr5y5TJod6MccGwZRB6dhsVs
NKP2gx1Y51UNTm6XVB6kawG8f4av4vxuqJJPAC7b39LhS7IwPxzxeveZs6pAvp+hlkZP7kPK8t1C
s97gF2hd/b6SUIefCbN/gYAOgZ9VP9z8jc2/nwP3Qi+CAj7Yh7j2s6ar/mFFaWGNGge/PHPOT1AH
RVMvPEP4OAKkXPEQMAHpOzBS1msEzYeRsk4utsuOBRuiD7r+aGHi6ua/cncC4J64ht2ZeuRM77FI
ZPuKeb6GUCl+gesG0hl3ItIUwE7b4KAhkFc/cnZwvdNbysv3VylWuNBAHWCoFzAQX0Rok5bYYXsd
ewrQsOOlM5ZuEUCsqaa5m4zXS3V5/W67PGu7zc1rH//qyhhafkdRJPjce/RFXQcx1P+TvesADKu1
34zlV4Rec6larmV8QyTKVsln5+FHLtQMVsvx2aOHKfUHAKbmpWh1fsdfJkmiGtCwEFbb0KeA4uaU
90lFqireCgyErjHvsdWDxWYC2tE0qpoVgG95tSHS5VygG0JgQq/Q2GIWKVwTEzv6P9NNVzb81HIQ
did22Nf4sPqrC9ujRsjZf9xFAcxfqMIL5/JVzLvskzNz8pgOpj71d6DIKSNJQuNdsfbEXNxxVUkx
kviVGmiXs4cOzqik5NmmKPCEhIS18t1MVpUhIRtTur7rFrbFJIPiLgQecPdy2nti8iAdvEFzztTd
fdc2lTT5WQe+fiGt3PDUnMNznEwuHJT4sJdf53gWwodw4nSDpT3msYpZg5/aFmQmG+0P2cO9oCk+
ZFGr9Vm1en/a5D+uYssk4wXDNQnIU5IXjLTlG6F9E69QKlXQsd58jKb/INdiLG3KQ0XcjHgT8IAE
llTg53ChlkfY6TbOnGhNAAng4wrKJTey/1O5ZpKjbDBW4H0942w/2WFVsgyexf3qU3U1ehRPKvfc
9TZY65raBfqEwdGUgCWG1NQH18FWDmNH7kIs0kwMyZL3WNGVD0wpGb8NQgRF3wZ9BEBe0uA2vo8d
r9zDSxQIZ2KyDo/DNSdhp2aXVw3UyIm91kuKhGm8GshLU3sqPkbiJKCoblKH9Nkvcm8M3p+njIZP
F27fIbEsUPCMFsfuF5mtnvYfHNwaBiEfOFrdI03GKaCSZNOPe06o1IGBj13DStdS9X/TBOWBArvd
mPkYjtCsaE7r3cz5d7yRbzjrNS291amLPwZMCz72QzQV8H3mb5tu6MrphbX6hOCKW6e1KYTeU1AV
pezDHS8ZEC3Fc+3eAgd6EUCWZPkXKpQfEDyShBvczV3/Bvqqs86/wIe77tKq1JMVaFEfrPa887Zf
KuP8lnOaJWzgokXN0FqeRvRiqCW9I4vBHn7lG7Z/9cTcg26eCTmuRYT9JNWDz67a577D3O5O1wBs
Dj/ocXZNHqaw+TdeokYzKCcFUrb5/MQ9VU1jnbiDW4RwPpDqk9r+SZnGN64gbdsncq8N3AMxqM41
V+6e6WdH2PDek0aVjTqKY0sZ71i5mdJW6KCwO5wyP70QkLRCwHYdn4q9yO7gWjdkC3pwCEaLFupl
0bQiL6aLf9YCTZLCjjk+FO+KOq7cprovYt2UBmdlqwojESJKemTSloiegS4Jzq6VbYnsnjcubro+
ftVt0Vkpb+9wGV6XdTHRdKmhg+VIS/bsQO2HeA2Zs2li0Ud8ljQDzhHZBrBJ6Tpl7JdOIF5F22pX
DLtnDP2lKgBO1NLn/9YpUHS4vDxPxFjPtVx5bQNHIlygDTFW3xcSkqxlhig6sW0UNLOFdy+eT6qy
F/7HNUBmD6id4nJNBXt7gzCf15t4dKB7c0RvEeWn28zur+OU3Gf9qfUZ5dMiGqJnb6n4Ybit09fw
hDdlC7+nGbvCTIIvG8NZ8yZGrzaoOuHHD94Gxe7F4n+oP11UtJwzZHD3xVBExwUioT8JwbDY2ptW
WcmRogy93nCpttX6xzrnQRM3fvKp4TQTNy/EOlYMsqX2M+Q8/ccdXtA8s9mcDYCNSm+4LzTYGTjQ
m2iDqwtFyofSvS4tmzHGFh5qRgq1necpK8gBz4figMsAksXMb7zMRtHeBGkGK4deKQUv83K4bI7Z
mZVIYzWA1V7rr+BqQhc6XqyT0pTwGU99T5b4ZTa2JtwG29NefyiF4MLw8Gi8iAOdKCsqw0DTSpZQ
OfbnRJXAwYsBwH4CtVGm7btXiwGa9IbNOO2vgQz0oxrPWnBDT5KjjX9paCsCSI3gsuBHbIZeiCAe
BbCLiicK9fUyucF6OIfDimWouk+pPynAwNcf4nw1mFaQh6PPtcm7s4n2+IdatsgwSWsPtTyliewe
BnYQGG25LTD4gJ1XzM+9u95cIi4RssfGLBNIthtO9rlkYChI3aSXtEdcwAAko9u19nP55ck/sjmc
DLRloQI44j5xG9EutTmD1vvIO+4ezHpELqinSDzT4oceAvb/VZZTe/2L5zhWs1Y+flsS1L0tvhUM
8KNEa7sMF8xpVRszgtc4HngAoYN3/BHSpsJ1hlnl/oRhjDIF/2ZuGZ7Ns1MgypjwrBqcK6UFYM4H
4XAJmRG3IJ+PFPoJuZzrDDL51sOo0JGmrWw7gsxPE1RLAH+77gsheicX/oaZhQ/mNHqbvWlID/9y
Qw5zrMqTcIiWRTnPjXg9yWzRdT/wrbLyVI7L4TnBYHP1SPIGfQlkS2gIZ00igyd7yDaTO3fbCw8/
OYwJ5HOS8p7GEEsuLX/JjhQuBA9b7pVGaf3pwQepK0nWS0Ybzj8jnI9EP1gYeUx8y97MkjV5HDBz
jThGHCBoTzQb/9cFUyZU11bZo+PMGWR5++qEXRHlM5syju7nfNQHt+Sa3hLl0V4OYHL82pj6Fhlg
lJutcipUAlfUaN9byVZ1dReAw2tar2UfQp/wHkJ1kjpMXafo2ptfRhoXBT6glE9W3IbnpgTS7KY+
JTYsHPls1uXv1ZW+0C2FaVijq/2siacsdVZ0lTbIjguto/1HNW7TxwnkV23TJp25+Nzk4uOmKWpv
Bm/M7UX7RFPDFJFBNgU56Vu8uaoqusxSz1FZVezIq0GNlpmbsz8PIFSX9CXm32yAMnh3LA2HOwaW
Fda3KEpgc/EBwjV2vQE35b2AESINWo55SUeAJmm0FVm2IThAYrmHEkFNHNVgyhRPu7WBrCLGygtf
vfrT5VtqZDYwve4IFVnwaWYpRBCQw0JOrX6YtYT4weusK+etGA8RoE206UfJuTWvArxQjotG6uaW
PxP55diIAE4IyQ/suPV8miz1DGBifhJYNgxWcyDH0JWT07cpwqqxgWLwCMvTPag32wgm80lDNHfm
lq8ONR5aIV3EDWSfTNh4Uyon/uFALT6F2PTFEYbmmtpREOUZaIHg/Wi20ZF67jZ66Hxt5vF8i95W
Voy1yo3IZJZrKWnvpEoaFdT7OFk3mbYut78N44nZqTA6S7we+5TRTCMQTTMkLCItqjWmjOFlX7+P
Hw3RVDbd9zuQyke+5rfkjR72lwuXBvPt6kA4Ru8VVX+v/fO0rPVZs44I7hlwToLCH3xNNAefK+Ys
6eN4JXP2UcI67j8RisT4pm5RXBvpNl/5BJsKiYnXzf8LaVj7o8D3GYRtUN2PJ7BiwgbbEIcDnTBJ
6tTJOkGk0yrtAHahB585hOn2ihq1zz1+eukAGdTYTJ+xjvk9MNCfsiDccKDDEzeZD+4jdlipKD8J
QDQ5Wly7z9Xoz4MyEI1jaB5mg1uP4w26ksypKMPFJydsWh7kfCMxoacvYJg652V/3VkMH/PuiFlC
cIIsducP8Z47VoNnxCHQGP7T5sycUMRGiRFx8Z7oxwlbq7tab0n7pIefSomKZmpc9toR1am3n0Zr
YiIdrhZZLSxbniNI0WWNRy69YC9/ahhvbMDIk+4svAB88isbSPXEPapb6KOh8Vql0oyquoQkU3o7
LhP2pyShstqDSg8O/W7Qf4ekLONiGXMXbW2stSIWZbkkVD0iaODL+o8kH/8E528PFJiic5GOvYTs
eLk85j/FD5/rtMEdpt1Nl4aVpb9YIiiafKcwFuNoe7amm8qAmyG4qkO189pCggiFGf2WiA8hLxMz
lQwRMA3xJnjkZ4J3OjXsK5+30R/h0bzIAUDZb5r2MMrcTjNexHCyzCVE+qxT9jrnQR2yXqpDfAEl
X+gEuaSKQ+eAQOhySWefPlldCFF9keUHKCgWcdoKZcS9pNSwcqOf6ZGRxrUayvnZKfSuJwRswlwz
sbQ0Eh0aHtoOrIQd78JfMwax2ZPE4Uooonsy+erd+Kb6R7dsv5wiLvupLgzKy8A8bjIzaI91SWtB
FOPAVBEemPsIiotCNJQf5C5lXOJGx3feJXV3cl3FeQ2XiO/JZ9216jYLH6wHKIPFLhhs7LVAZRYh
EA3Vn2xuyzBH43vQqDM24/Gw78jq3vwGqMachtD7tDjNOyCbj4iwBuKOsoHy9pIU1AFeYMM2vD9j
jS4xJN//vpm0Dv0hi9bZObuJ7Evt97tkzTNqvPiyCE62hZuHHCgN5Cp18QBfRBlC0QQn50pNbo69
qoeOGiUNiUP1DDXcf0+Qz94DI/wo9z3sId3d3RrerHph0iy6wStjCh3Dimiw9qAv4BmO2SBjb9Jn
g6haw+/WCdkvS39yDpPywnbp4QpgNoqpBqerzBaVJPzOoxcPvAuaPQI/jd11jiEvDiLhJ9ojTYn3
Cp+zrXyp2uK3kZWhhPbYHDmmm1nEhW9cCUBzsBYC4sOZedUaNhXYZI+NTeg7nJAh98/F9LEWXvtn
XTdal/9IVfIf4dQa8JIXYX2HT7cjYkyK8TQMEKjx3x+xLb9Unm7wBMnInRgpbS/NQW/7ZJ2qeByC
sU4pZgLlcJuhY0+pK6HBv9Vfw+vQxmCcI2RVLr/auO3yIog9BmCntKhC3TYFnBT8gRxvRyr7AadY
ZWLFueIdhgSxHVJv9j6qT+b8RJTQrpKyQsmhHFI1s0N888FQ98jOuEWyzM0pQtjRj5z5/NtY7EA/
YU730qKuQTJGvwA4NGr0gpy+oyBiz6LZ+0B6D1ulafFzZHFDz28ZQUhl2KY4c0pzixMifkvSp4ol
ifibym/Gi5NzZyG8eMVDsOZfbP9C7S9fca8KrqK00R7iFNI4YZK7okQlwet0da2hItesg1ElUNos
L/S3dTnm6x8SSWnL6hGVIUgUOC61b34WItar13mLSRLYS+sfz+9EDxtWnzp2W/et2Sdk9exHcJwh
gkhCyNRqLFRLpCijwT8oUYyRtiEDyThyMorjrYCO6SBSbkBaIeQK8MZGnba6i/Nont39Cz2hIVXX
Q38oo8pQ03t9c/eIV5ZDotsrwLaIxfDUWYj33gEumldi4mneCIeVJVFECHTH4hMbh4kxT7bz2zVi
mlp3awkdXc/VGfV/ry8BG5QsPGOGx4G1asPaL3pKjX8ODmiuOTLLgef6a9XS4AcUv4avaG3J/fM7
TIx7poBhu5UZkfIlCtUDh9YuRlXNlSFYATegolJkvlLgT93FI+AADxdbOjiBQNMDcRK+EO+cYQ/z
pISecPKHjhxyPfFsfSdq6mv1YsJJkf5zKUNVTKTq3I+fWh+0wq2sxbPFM/7zW7FVXYhQxw8FXrwo
N0wKwwoouYIJBzSKzgxtfRQdPLkOrcoCfbDnXO0XlniBwbsPEy2Pgfqk7vfn0YI6NGVZ8Y1CNWaT
wDhCKzUyQ/Uy+gYhKBbWgtdkZ8q0LgeylPvjTdif8tANPsCCgqPQ2zDU/RjoBdYvCIkPyCZ58FMy
TdEp340vRVJ+VCqQbJgmW2UMY6Vj2vsRh4F926bsGblqNOj3m0DawliHXweqa6V93U0WIDTtxdnt
06QWegrqoFzuP9CGAPOfBiqDF7plccZIBzxWC1Sj+4wfKWNLfGGJZSFsMUmpxJKB/R+Gmt4p+WPz
qwZ4x2Dhx9mdOuI3UPVNs71pKvzoijns8FGDeiuCy8+ScCZjJF4skPDyCeRTZv3i0PWqcwqGWiC9
KE7cq345JRyeDNipLr0GuttrunX08bAWERyJbLTSwsLuBo++0uf+1eOsjHy/IHPl3Mv4hypLg93A
qHyG/hH2ftAyKax5W5YLYkCuQnPXhoiowdY0w2oESgJzN7i7tV8GsYER6SVVR5sQIN1yrW5oyG1Y
6+u2LnK6YpcX5Xp6X5QXzxv6ILDkkYDdx4VjgKAqIdlZ2SfAf+i8uzXEFuDYF0I7N0aoV2/4slS6
deAmUqgkaU0Ib1zkzmOW6dlqfd0KJM0C8q/9w4HaxwKELTlMgAyUvgayZfbMBmIpMpQvX0DXArzj
NJQq3xKdZzA3pyAcZnDik1Wf9urKjml+yAaT1KMsAo3xGr3CNH2c6wbo4Fqo7OHueHu5xRZZhIay
IrkrAo4u++NcDmsxcaQDi5E/uBAAsmb8JDQeWIaiWogv3b5F2FNeurvnd0U1ZBOgGEtfJdOLIt2G
Pk3YskBFS8biPcZUHJFY3gPRen0Mz0JeHbwWCMgOrqghN1b+/SASxJHakAHO/ldB0iaIv9NscgXo
+U0KvyevCpMxy1XyjgNLhByVNsDja7xgAkqoHl5b64hHx/6q8156uo5Z7YyAxqlcNseTNtplMQsQ
KdBhV805FWAqUedbDnOvM2WmPNENn6AqxMr7WLZxF0mEWEIKfjRI9Tih/MPXmUKrojKasnYjkfw1
OxXkQq2yGepXq21N3VaIspLGjIiVvQDemZFh2AvNokd6izckz02oK97Prp26MPl2KBG/BKVkSkqh
LFEv0x2VTICzC99BYMmLuwDyUCe1DiaBq0lhlrehQGD6qIOUR8aBpTEUbgv11PFaohEBDMAzQnB2
Q3pTqPrhxe3W90+XUiJrF2IbLokMxHbs4MUMfWBYs3wCAt0M0jeDN81yuwjY2K85jyCsIaAHl4FH
+j/45fDmW22LBvEV9QcDJvoQt5th7D/Gh+onq3AcShBsZeEmVOlYxdxC4Oq0Jvga2jLpqj72o/3o
IKgGJ5u7Kug9kJeSILtfz05AGFaX9Yw7dBH5b3FkOGTVd4Bt+o+37EWKFmFBxbSG2ulEcjZJ8LV5
dXw4y3F+T0kUK2JqFcKlMXleAVMXb7wd/o0q+bgRsUUViqrdEbV4bsPPxz9TZNzqVXo+kSySuA9e
DwctqFa/+/wiIkBm50HCOBj3wlZOAqpjqfh314eScjUy6yzArmc4uEl4nsxMs8x95kvHsQDVxJ3o
/vpoACVmSM5v3kMGKCdjWuJc3AJIHK/VdKkicIYE8c5KRYS/Bp3Tv3pXA2Z3fAVdbheursG9grhz
tzKRTpmfcTTJGg1p+E2VCuacuZCRm2zUaq7h8WNpRA6LikC3MlskdvPWo3yglclEfLwhL63FP3yk
XcW4z3MNE5dQF4PhNqkttml8fQ9qksKuai19TeuotusLHEnAJBnJq0QhWll4CmV0+W1owpz3LzYn
5oC7VqiWypnY3no/uS+wh2YTc5ZxQhX/Y0fgsQm8/r5P1YtDHSGR7JH8fTdNXCzIDLgGRAkdcKIK
E+KihQUFaWANWK7tOZ1DcYUjPgvC0ukOhEB330iNqF1JMFxfIyNEha42+oj35uNI1bRQ0uqq3zNe
Np5EfhqAB0y3fDbvI4CAVWaK9DsVl1q+TD8QICoNZNWW54t4gUzqOFdIc465ANGucAmpt5YkpZGa
uNTdsHdmvTDFSgW6lzuArydn+FdUMIdVtEXnanrRMKz7hXCnXLGo5ntYfyYVVjJz6sKggGMyZ0Vr
5RupuanRNKh+RPB+fMG9FTjuy6VJ60BTDXttHaUpL4Rc6fjD5pUfmfc6b04k6//FmwHhUtBslHiN
TAKGo51jrmRnMA8PD7gQRWzlo1VweRO673+/nVPkZqM2iLwMI3TgsZUm5xnma9T3da8rFL4ZrYWB
HTWmm/I46v4FN6AsqZT2Vn8c/Wj1fGGbOZm6g9xxq8Zqr3Pf2lYxMLHuM0ap66w4Mn5SpFPl9ib1
E5PtOrd1/wBGRWXaH5fFgffAdeQyx4/fx3mt5RQeeLlPrmEjAs6BpJ6Mt4oFD5mL2sue49rKPjay
LqyXYk8PAVcethdsc7Wv6I0+xgg3bGwMk/NX6n6K3fjhZdOEO463X6LAdy/VHSwVfPtV9ncR7MFb
dvdDTCubCt58AZFZzHSZrsj4EY7StfgndXxYLMocP5EMRIgIyWKkbJgG0MZOOd1TPpWLpou9q7EJ
VGCRrgmFz5mq7lyXSA6xA1l0qjDrUqsJTzfzJ2vmBjfcgCYmaXxBn2e606M8WE24tYYhuntBPb6z
cYDmF+Kz6BB8mfi+LzBCJGQs6rf58SoAs0+J/yA5tkxbAUcvmIueHuBehzByU15hDAgf4sc1/yAj
0ul1zilKkUYRvVdlh5DqE+imeXXqZ3xCTBErKRq58ktyIg/ojPNzAVW3fmwFQkusbyrjDiRoilQ0
YuVZc0TKcJ3eAw4fVxs8M6C0R/lvr61jwWZKT4CKsYA2nTo5Dgu41exVCPYx7RUE5aLjQzbBw+WT
5b69g3bgRE2UVJLR7ylvZrkJQwA8xiLEC2Z7hjl1MImYvCDxz5VV7S04memsBbRFFwmTdwkvBTAr
XQQeKhAWTttmp5r5qgHqS9f+H6Aar0c0PB380JGvmkqS0UCjUT5LEYBF500JdvRmPNku1cSokcXF
Q+0dOLlzMgX6oRJOyTB04cpRU2Bz7HK0ii/HIJyvQdxozIiKGAHGu1pnhWab3TOVCCYhuUWztj5u
Ae5qmE+dfnnmYZWAEyXFB5r+aDMq+QRK8Z2fCjWgqf2PUj9nUmbxQqTz+Fn0LTgwJeiEiQE3Rwpa
WQzoSgoc+7c9PhUhXh+Oy+Ht5jmvdWCea2NFkQciyaZmaxMJPdTHf3n2O7MOXmQTqdWf6G/qkDTA
NKdt9Ix/pZKpvSrNPFr5fedyG+XnZ2opWX57LweNj5mB1fEROAhSWrTZiF5m1YzaOXtrpHmQt1zD
ROCDA4QoS3L2qbBBo2qdzHlUGy6ZdKuzK1FrRUKnLntvdAaOgJZU+wv52OabyicdZ4XnzLi1p1EA
LZc2FJ7vSrkJ1IRyaAUhlZrQxBMWlOCeVaKIww9LNbzOTvruwli8v2K5ckn/WIzEwbJbjcdczL5Q
iIDrwYGMPS27vUNO1dT2L4/VLnZdwm/mOw95rRU4z7ilP3kwQKd2EpF0XemPHKvk0IHxbMjzSzAU
7BK7tI/nAfKKDu09HjtDGEwbVypxxZoEgI+6C+CzytGBfjbMBffR7mdXC8Ie6Q3dwgADW3mQKsNA
AbtUFuT+V1O5YX74sQvCXSctAyiXCTl8dcWJtcxVcZQRIdcFCCNfnwivMaD7NY2neu3C/KLjKs3g
Oodn+O0nE8lpZxhkyK8OTjQDst6UHzftBJz1kD5a9txHFuvkojUEda9/PIm4/3NqUoFJcD+NAdMm
YgyLGwM9zl03lPKHvujRMMQApF3v67aQo+y+NEthFyf1uBrcwnTCAanF+CijG4eM04RExSJglxcv
B7amsDCImQ5siYpFlxQWp0gF81TtIaoqc0VWUPBh3ugrTqnQ8dhvzVG7pVJ/0B5drr3EgHf00D+E
M+RQChJzxpxsoRwtof9Ad2k5vWrsXpQGQNtO5Yfxd4xI/v43ImN3q8coSTB2rmNc9L9D/Pj1nRkt
5vYl1TNCM5YWBnbuaba52YZ2ixu/gI+Q41zo7m6YwbzIXvmkB+CcS9QDRPNNEAdoqaHJtIwV+ouv
C+USKrxKE8kLeEdcqkZU9LTXS/werQDvGFxoEh563zGTdNJBGhX7cXgaR/Vay+TbL23q1fPmI/Zj
ugQ+YoWdlKoYyhnQLCqdMWhGM31vJGxJWJc3PPEAqwTJUBgzYH71qb1ySfZQP9elFf20hF0jPuE0
W8esmYsc1QEO3B5bn4ACg+4IHZ2BMo2rsTvaPeK/GPbIJa33mO/sO/tgbexay+iIoVr4+gFGCC3D
uZDUMxEh1n2KsJzEob7tvrUpE7Bks0MJ548W03DZvSJpouKdmcgbrmhekPWQ2LoALfiba7p2icFc
waWaljDa0y8KPdKX3OD+lha6++/upZcb72r7p8PNcIkq/5I3mG8Li/VRDk/3AgxWctoze5EqPnVR
51zPOyLi5iNzAidrU9tRcgf7B5tVsvBl3ms9gMfdrcKSznpriudxHfyA4hxoyTfQ2FYlPJK24Uq2
Tm7kIfCBR/3+ur+dZ4L7HZXCWiHGJWX4bja3erI9z7/gxm5vHaA3hV1FOBq2HqX9+0xbbU5R5QZp
676muUH8iIlo2otRUvCM6UcrZv4ahCs4pw52LipuQ/vC8x+inmVSZcYabl8h/xBoRA0K5ncOse4b
/l13O+9EMDqZ4+SRvLb/zyC9BiBxFyDQRSfSnF8dJ2P28+GU3TGbdxgBwH+igwD5yahgUm2qxOIY
u6gdiNsAapFrciiPvnLcBbkbLWcef1lzN9qvSBywkzplSI+/su6mUMeJSXnRL0DEonKzPswzvseg
1vDFfOhB739AcsBw0cx5vYaVbuDqM5mJIlmA8Kqh50X4SC+e59qycLGoXtvzXDASEXkY/euctR8J
PDecQaivX06i8KAi0HeFYOFDBmVgy5NwdO/taJ+GE+D+SwoCdB4PRQ0rPMiZxgWI7WVRZ9Ol14YP
hrZcHQ5yrCSt8NFtf5T8GPdrreJWFm06uNBlx6FsvxtjL1B6BY+AOboWB6/mcOKw8eF7IhCE5Bn6
9k5JyzV+rVlbfslQDwX9gz/plmjARBrdrOA8KLCLVHsRaEveM1HCanKoutX8D5LebX+2eK4BluWh
nVjogjA3Lrl49J2G9oziGzeqsNLiHXcARKep8HUXEyWfRMIT/ToBn3vk4ox2s7NlSfzhi2Gh5pzc
9DUdA48FizLOsa2Fqkg1NSDpVXaaaxt3LWGqN6yBFjcbU2BzZ/XugYxepcl39liJfHfErUaNthST
hiTO0s27gLyWEfrkkm95Fj8rJKOgwSJnqZDl5Ab5k8VbXHm+LCKl6ooXd20XPB8lQlekjkSt/89M
IO5RFu+A6Vn64Ngq843OijBxXTnY+P3o7//0PT1ymDTMQSL0+5kx34n6f0FFrCe/3lGzH+cFecyC
ehjFPv2zw+b9D0CHrfm1Z6zAFjl+khMNuVkA/iZQ9lOT8kaerRk+YO1SaPk7CCMtcqbXneWa8ctY
aEu5XBwBl+NqwlYTdiJnqz00sIvkLaio/GuPb1c1wppTFumJYLmemiURDucgg65/cnd0239i2/+X
g5rP1vdB3PKCql5EMg8ndDeP0iVTE7Dr/uPRX+WBUvp5xSH+0vTJ2FXBbSJ0Cq+iWbSL1rEZdErC
FrARIkIiA3cBJbo2pPuhK7eCbZM5HT7n/6Up4Soy/6dHf1tdoucDMgAnWS211rD4RddmwxHvf8T4
d7o56WJrgoPPBetHaFSH3xmuzr63UhIWKYPqTcIttjhqBlETv3GqzeTBMXLxc0j542JfffFLnAW4
QOZ1KlU9V2zmAHxER/3LfwW3g/DqntMDRzy6V9qc6NnbC1Zpezz1jrg5MfUfI7DspGj7ZvV2Haix
FKTor13PGW659sapW+8B8z01c12CIh/7gYTPOCnzgyJ+IK+MIWiaporZ0x1Yk8cXg0CCqLQwvVju
WNXmqvqyAUJO6+Iw4voyeQ/VG6p0p44DTpGw4IRa91MFiGPHQNelwfQWlyaw9nRS1d/jajFw3Xmi
TpljmnF5TIgpB41AFkCg4tnn0JMbMwHb6hJicPjQZ9q02vjyE4Cn5eWmWkBRT6W++PKKwad8P5/I
qOXcWWq67eoHvhYoHQCsdTeGwYZwJkEtxrgCytNEt4Hu05UxCgz8Zcgp2PxgPCjV642Vi5fhXjG2
iDe2sy0HYUY05HKHJQwQ1/RXGksL1fUmybK2Peskx1sfQfahzxPCbmfbfyv3mD+P0FuDl3TXUkBo
c8LOWxTVVrjepx+tIddORPz2IFWp1PN04TtFhqmaMFu44axPXxMwvwZ8Oq2kFDev1s4wucI1I6+d
90K3T/HFmMdUFCTIAFixhmCTvkXykAYfBb4pxsIHAJi2qmhdvcjblfZTYbFdYDlFJef9pXiptTYw
C+TTASBd/mJ3bCE8aijA13+sDciXzxUFaY+1cfqrxABD6e14SMB/it1DwKZpX4SQX8+VqUBj8EaV
r1OFa8O1ILI+syw+mU8TiQ06EKsCnYhMb99idcb7GmcC/xOfpZXxxro9t7lyPBWIa+juNhEbd0xS
23NmRgdXvRgNPZcErPOzrgy3x3xylrbsBmhAmDfdEqpvILDegK8NqlzuK3elrFFiVJtrbKO0uya3
BN5k9ShzkWH10Jz/FdINQ5VUZjx0fId+bJ6E5gfO92MEOJzzBUnT+yjSal+7R/iEYzUkKmeSaCqS
HxvXOtiz53JvDmQ/l0a9u/Mrt+LYmPPKedJ5yPTTWr7Re3bqkL2fKswNxtadUwulHFcak1ToW7bs
2TViT7mPvFkDYwfLWVbNSkAHgzGEcwdLPucIeyv9nXghfAaCunA71TtEajhXT/4zwDswEizDoxtk
/oclSzkQvJPEx4MKq/Iqsc0U7ddPwr4EyYRXsNls6aXlx81qqMA7xiO+S8lbpvsKwsVFFGwubr2r
THtpNLkXrFSuacmr8l6Ick9+8Pgt8bFlXgwigRvlLxLwMLuXwM+Bzu38dQVfUbz9D/Yvb9VmsbJG
CQDHCxX1XkmCZnNAk+POQKb8PrtDZ0zbt9S/747BEi0uN7Ev+0aIy+49khmsLixnS9Sryj0Uoyke
SCIFPV13EmeCqq5hwmhIjTiKDf8EUfNXgmgcf1Xma/eD/Q+fKAULSUrks5sRnHUiG7zC2/yCRfqB
We3sv6+jFFNMkys9T446jD8qwPPAo5mlrxWwDGVkD9v8WYie9UOmknwKQg8hP9K2wW63HGBrjWsY
F0auvrUWUkBVhQWLwE1JZ9ABdq9aCVEyr7XLwPZiHtnurAEdi1LvbxO2dgqnuRro+V0g19A78u/7
9xHuOoAT4h6QmB4tOcQ+un7SE9JeWJixxbWhub90R5xsuEDKWFPG33eltYyL+5Gcb1Nac3JymMNO
/spMBLG/D6IpYiFcmIfeksxvJLVnbxP8H9BfXNH2K4f+t3XgBArCoqVzruAZtpE8Q37Tg9HYDzM1
cjszRpYwL406lt9AXBxuldQ92uN2LIQhC88Fl+aFg+Uq0w3K044IrFSx2aATTNxDGRSx+qz9vc21
7nqqXUH9Kc7ofpCFKF78wCVeIZPBYPQaQd+Oa/6BXBADEumsb4bFEiRqbDIrl+Pq/Bkpd0CMNXCX
d+g0mLfQFqtw2fQuCuYy/N2ZGzANMLLMYRKfs46gX1K8+3jTh0qNltBxSe009ff+LxWI9WDIrCTu
+klsrEpe0U4pux1F5JTwwwy5WWo3OVBULpm8VUtPKwnt9YpX6RUq0VJfsEs30XcniEwqRkwJU5PK
vV/1vP5kMLb99PSn6VNls2Vuj1onrqRwnPi06taFScj5QuhteJYpFji3TUlRCTztKKeIT/kv9kD3
m/FyXM4NX0eRLICnW8ZSna97yKWAUVqnV4XrT9fKAMXdzs45IxouTCLOrOB+NB7nc6cInRunILqw
WbbCzS8GCq0I3cNrLNq1b1jEDfEs4GZ8GjJZWMjvTTe0fXAQpAL3hl27O5JHzj8XHPpZHc+AZAob
UZF7UJQadN1UbAjyEzh2UdMMer+LnCo32/71FLy4t8nQORY9QyxRY7+1KlspWUD69jyHOCVHmJ3x
N12KSbP7ykqx4lF/bJzFG3PIxvUgeOHSpY64ftTmhXB5E2g0ONimpo6wOuraJ4a6wDJjEXn/+fra
Z11tHEw9AUz3T7h2YtuZuZGGYTFuKBSuXGLjJIs39i/K0IdTVQOorPWOKo5HMnKREZzKieAfEw1n
rtXW7J88vtLhVLi9S4UdzrNUWxZl8nFOFBMe+fZ5QvNf5rH28/W8VLTB8vP3Fz3/ri7QGKlzvkVI
MMfvFCU/FJQQ+D8HWu+6ysybPuiobU1AnIqBqc6G3r/h/aGk4wXnWkH90K/UO5DtmjgTlMPW3oD9
pPhmsBEgmizlxS3sn3e82VZ76alJuqLp0rFnnocnrnGndpX9wskX1uNAFAoMKW5sOBBsrVvO3X4J
YfMXQTty5J0h4QWb50i/3tF68ZvuaRWWSvRECpxmdLbGybV4QzfC1hNDyaRQZrsr8s7nGHOVr4kM
wBZw9H42gaJEcF0z1O9WCnZq5074ORSbIbRTRSfdQk8i7jWKBrkRcNcbzxmXCz2MBPmBIDmFVL1I
alAfpQ7Sffas+3UIarI9TlHLKo0bn829jDSwDJVBNGOfrx6hNci6XIY6SLaWa13mzY1fJOTTkVfv
w5NyLHvp3BxLGInj6GamxYphcX0IX/1LjBD/M7pryrx5EYMK5ARAqG2+kQQ6AgtaevkInbFqA1gt
9lZrOujhYoBmx9CjlrteI0/sYbpVguMDIOs4lwlm2NTBkGhZPOir0U6G9KPv+ehJQYXD7Lk9sN6b
aaP/TQJ9uColNTN1C0/+jHRjSJ1+Tes/eHzs5dm5y4lXZoB4G4xC7RPsICH0QZw52AOXsHCSjBAB
Ox4Ac9/CGQiFzdtKkMzJMpPMaUxl1tqBTzMxUSQOU0Jxfi0jXA9CboPWo+vnOXKUZuEevsDGx9at
OO0Go9QAJ/Tuo0wZBP4lyVCl1MzD8f9hb7vjQBEcakY2afoMCLrOjrBgpO3j/jSvkO/lOMi/9WJH
KSp3BA8/pigmiaBMj0PBafnCYxtcpKs53PzspGycF5fLlGoz8tNnPQIlWE+yroUTmqQ+yHxqim/j
HbR1Nvt4XZsRFuYDlity+/WzQa3C64NNNlvpU+tPCp99F5xdbU1Sf+vlh2x+Mkb47oHVEogwmg7b
NZatvT+UDUjIDoiuVj99Vhc5ujrroAiHS3aWbJvSnq40JeXR4wE48KXFpeSVVchPXWgpDfzyb+Ex
WFBs/DI/BhTWAPOKcILZy9CnnTHSfIToUkde/2MwN1fRJGTz5CDnaEnAv4IaPB0TxygalTJvnkmy
0nCQ4rPIs39E56cvaKZkRGh7uOmNG99HorPUHAlFAse9eO5FflZhuFH07B9GDaIOYdEnuTTagIVi
uzdNDSGEPaOxeYxx571xO9Z1o/QRCNfyl2dOM+caC2BrQvA1E0JeTAJI8paMOwgMqxHYT3b1Ok6/
vCNFcwaIwlSfw3KY/cslBIU470jh+ppBmC0DVToAVoZ1aR775Bw2+zQt1er4donK75L6yiqrLeqf
7UXACzK71korkI3BHRoIAIva1lv+2/QgEcjgmcz/eTV20M6iH/WO83H1ZUci7bwPMwGkzCyyu2hF
ew9R8Ath2Rtlh2Wbtj+fiJajmmp/7Cb0+vB8LJPZfOL5BETrXUNZcTdq9f4RArAG0u/l3E32GTkZ
+uVa5H4v3yAxknIwMZ1hDnlDwcAMj3jmYAvP/91Fl5C6ISvqsxTDp2XCzixIxzxIjWjar1Zzyaa6
4VaT+e6yAGZBNVdFOjPRnltv8GyTtszKcwXX1aoasV73UHTcAGcZNNm2oxqA8rw0MafgwaezlVdQ
Pm62bBnO3wesGPc7DezWNF+mOLmUpbejdzQQw5yBM84OVP1WGhN+lnDhqYe+prncZeMVLkPHrd3V
IITxCzHcAdNEAuMA/u2jydFAVQmZGwD/WDWcc9Uxf4zv/gFydM6Isjvl0gK/zE1uBJ3WMxxmlP+w
EsS66gcuIjbCGc6J4hd13NQO12Dk6Su7Bo2mPHPrijy9KVcCLdRTHaU0JP6CIEjEbm15sR867PCM
BmUl+/rTmrWAoLK/EXEtimrRFmzzxk2gXl3Rf9qra/eFY7Ha+PoDG1DXnUXbBo3IES4SE5JnXESI
7tLXYfgvOzGUVCs/khAZrWQrkyKrZK5bVgLX78pEp8OWP0TqIsxWtV9LupArVhFTYOgxY1QjG17b
1PX/fXZz3e4k2dxm0adS5S9kNXUvnJn0alSQt2dtpEQ9PqHY5A8Dy5lcctvQ8K8V2QRYf/USlpMh
bysD0QTxE7G6OQkhB7MmLDor2nPriOA+XpWjEmR4SSSTBapQ5VLg6EAnmR6xAm3nuDubJxHb+B/r
qFn/RER2EHS08r/8Blvf2DtmDKKEIOzAqyOhdwLpZqaZsq/bdjgtuGibeXDr+CfCsbO+6cdUAeyI
jY7J/d4T8zAd6ccNox3azF+xoDr2CUFfY/YlfHPdJaQqIJ+Od7p5FShATK3joVVNSI6Ik0r3i8xG
S1wLLqhuD0KkBu8TWFU7tzZZXiP5tiusHf5uIPHtHAsWUnP2g1VNOM+UVJKxDYFTHzQ4NzUo/1Qz
AIhnCVOOMIs+urhyK0F6uvjS0hGf4GfXBMHLRilCm4vQxYJYIvKC8smQs4Jk6TsmnIrQv5p4Pmnj
P1IRykZz8KEBQHTJQrqohEB02TzmgZ3lxjmid2kKjee9RPOl5cY9iL70A7YfK0SBPTquAkiO/hjp
qUEoqgB7FvBqb2ujQkJsGWaTy7TgyCP1GeiCy0BQLaro6vumFbypmUwu1olPmxvUbsXtNKVZ/H0A
sZfL8HL/TTfYn6Ra0VY4ptZwroHEDuYSUf/V8w6OFZCthDmBjWMIKH4H5KCAO7XVpQXBtiPTYRdC
Hfp7n6PcXti8hZ3iC4uWiEvDgJioxRmIN8RkxO4piURsc9PfbfQW1umKwkob6qchYfGxRm8IclFz
CAORA6UBfqWGyH219JQf0mjqY5PXB8Q77oqAaTYbEd2CwiYJDuyd5xsXKdqDYGkEE/2xPXPBx7TX
e7Znw2lYAh6bnL1JrigbLB5sghz7Q6xKVir5YV2A6/gFnDHIU87W4TTjkZf/ogZP3y4OnIi4EhOK
vSc09d+fnIVxpggM7N0pHq0V7PHCNDDmai66KKf+0+6GgNIE10RYoyZUJ08o/fK0LscrVttEmf+J
w9DLoXIHUZ29+P/hKeulXwy7i0Evm2FlWF2iSEwlCj/XPWqhl1MPcKoYKG/DdTFtJiZoU7INv+Oh
jxwBcAPXomCaLbTfOkBtikZa6oIIU20qZ3FALlZzLbQJKRpTnjYoYtW3wgmuQF7sIis8AVHMJ7N5
haM7b+9ZD42P1m2w7Gax2b1yJO/TQGzGCwk07Q4O1mNlevUA4MOOpZuRrdeYUzFpoJo539KTvknT
TqqwHBQ1hebj2svjZx62XLAlTmHbLTkG9gzkPVaPIEwXj/JWdE2bnpdvJAlbyKYfNrrB1r1YG5ZZ
JrDH781wKRNmGRZjq8FbO/xKN+MftyCo4nE+BS/PpsjYdDPuZi1nBIBeVnlpYsKOTrHoGC9BAzQj
KONGI3tW1UQw+NicxcVoLEpBuurq87zA6VAob07yeQaX5OALLmAkDaiEZP0feDYTFhe+u2YGMCK4
g7Qgjr9u+OLtmHB9bswRSJt1VulLmHnExoO6eVeqKNFYb3Kc8XT76JndjYW19Mc++O6h9Nhu1KoT
yBZTW34qNqt1V2JXzBW/dTvZXyqDXwdaR9Uhttn9YOzdJMwJ2OyxqB3KbOe1wRUVJZY49pB5cd2H
YDxkUphhVS3OfqsHb6W+sYpgeD7zmKFEMrmp3ccfrcdTCjhfHn7DBU4O+C0+BkcD+HPvKDl0Es9A
RZIBceP8WR1TEYs+1Pva9vS/YnV2FBeQlOBmUmgfIrFfCh2zxsmjfCR8VRGM5WHfLicNn3ZXLL8M
FA08U0gJnneDBAW7ylIH7rp1yJXE0EHw+F5XlIYI+EaYg6b//sl3dXvTWSa1M1MhIw/g8jTF90vL
3WqNlX/2Z7YWyHfZUQtPBM2xSnmyUPlOyrn/GrgmgQ+3oniAclaAxoUrC941UquIua6YMMJHB+X+
FMrRAWqQv8z6Xu2iSbPoIrnlNAb88PU5ZkzTWEOmBtGjoQRRfiTjaCy5lMB+b6q8ytwUYIWYRpsp
NJ9oUllbESm1hGEhbpar21+CfXWnVJ9g/0pQNAQKWZmVsRKl5DheuvS7tjjuAJPmFXGfc1Hl9o3L
oMEmhI0PcjHYREQIY+OLaxwuBWXgEi98RdEKXIL29CYcy6Shm8VKe0/rpIuRqv2543ULKLg5kADf
QDDbNrG/tTHMM1nroRkPLiADMx7eyMH6JQgWkXN4ijeVsDNR8LVKEePhiy+TaRRGDny64yTUnD3y
SufgoBLNH+wRDtSkqvBGS14OPoQv8fYbHdCcsgDDaorCRtnXlr1FmTerxfGIBnc6fK1fVoeKfIT6
9+vh1XlcHxjuY1CVyGgyVhI8R2S50WAajv4hvug5VrUpFZx5WFte9km0/UNSrWyhXguOZ0eqzu2p
c7vI+vPGTLe1JYvpfW6Fx8vE+wMsfh9pAZDcXSlfUL2nKwOgE230L4JOvYDByytUab3V9KQOIxG7
xV0xfUzOWA85UeM/pYyn+Pu/AoUK4ObPD68uo0EQm6XldqtaUg00naHQF4YYYeWOT/lLo40LXTvG
IH6wQyjvcM1JucM2adholOEBI80PYtMgOppGZveHFvv1KMY5TINP0KM82o0ccsrPcE7MGn9+aFty
AVzrOtQ5xwE01OExkkX8jecRdlzDVQW/krMB3vCQgq72Drbl/021o0z711sMvp0uKCOgaQ3+sGL4
jPdNPht93+Tg2Ym4Cfh1lhJUevpAz2YZQTm1XJG5RuEHw1BT2g66ia8HmRVHuz843HBeZqUAUeTo
IZsgBT8RmcyojvVzzI+lKHnV1LY4anOHsaaIkE7RfCQBAszEMxxA+kz1RPBp/FMCCQV8iILpXvTX
07v/HMHgsqlVFX7CRDD/1LKb+FQLJWJSajXDtj+PdYZYhpRkcRUtG2OENOF+cTcqiJAVqnnGoDwY
/r5Q3q4caG0HtmldWgSdnBskEWsfV/m+iFvuFq4Q0vthuZeRgG4ePsEl/9RBKDF7yqE1B2SPntqZ
dniGC861Oe7rG+4W1GALU9bU46X1LaEzJa9kfcFt/0MEhrch/v4CWvi4wVDd6k8X/ygzp1+spAC1
EE8SWD35vUMgLtYnwP/5W0mzjK96gIsQiWzrWx4fOQ8v/PVixSI4z/wJkzZ/dDDDE+lyvwEbp9SE
jRjPCC1weJVnxA+H8FRtotAW62OroE9ehEZxhc81eGl2QYODmQMBYMUUVd7U6B77md/K8qh+f0Vr
twdMre3aC8EQRVsLFAaU8RdMF+FNCzXa4ZOOSRg93YbqdfQi5PEPY+UdSr/FurdZ2xcQlUYop157
GgD3g1yWGRIiL2IeHkNT2XD+F5pwrjkrx2pXvirz3XPjWczB80DpPnxVAtos2w08UUVhM+B2RF+K
kqUJOH0DMSbjtU5gLo4K5D4i7Gc78HmdSw4h89f0Cmw1o5pOcr3XhGqDgIg7b8be7JCM4ZvTJBjY
y+lpO1maAC6PXqNPgQA9fioE3SATeerWXryeuoxIO2tkOiTSbWjNq8C4IVahtbgBXKW+ewTnMzfE
4CNXCQTz3A1Tdibb6HXY4B4mqoUYg0j9RbS13XDV5uyM/Ekifc+0l+Znc72ycfgDttGT43v1c63z
QymbWxHpCApxppjzgR9PQa9MrJbN39xDzAoMM2nEC0HTTRPIUnoY85ue9MijZzmtYZ7gOhYW4kXz
rpo8gryx3SELxKy3ISxJ+uE4q25QMr57ujS/EDUJzqgBWJQIMRUdjY98CwUzsOziTsNHmVEjF8mA
SOEIZpXzlARq/AoodShmHxEvnAsz89H5RXr2pklJH6STEbDW6H4lSg3oPNpDlSQwM71fVohY/yLJ
Rfm3Va8t0O9dJ5fsJ3FVzDbxBMGBTixVa7OPQWLSvMiggwsQ0Ej5lzMl9nhR91lT57l2pwmdt3lV
Oo4OxElZDd7cuOzUlGXE6/C1vsptXKMhrHkep0+j0foPNQ9hsFO7BkJAl2iM7ZP+NhJ12GBEDS4D
oAX/yirCf+77C9leU9Vp6vgPeeIbcXYIJvstdoKRrlYocnaFsJ0KXPV36GQ4Hil65Jx5SPRyb5Yt
Oms0ygs6jJid0cOcWXlr4YymqS0jlhguatF8/P8gsxUh4qNtJsWkeeTdYTmpTCdp2RIHJG+47l36
YgZDu4FV9sGJvsq+ZT1GW9KX1/VZ/hYeQHRwlHnpaFMWj7d55h/DiCNKrUW9w4a6Vjt61kPOHP+v
roZ9bKhh+mBPTsOXd6OEiXViUe27LxjfRt6KfMKlwIBCnW+n8H4ifwk7orh8YTYS5lKJ7UT3/KrG
U/X5erjZZ54iWrQUAbmzDGFwL5sutWMcJj8uklzAxO/eH+R4xJUu2Mka61PcZ7yif6Vyv5zCxJ3+
H4RoG8eNL91GQZtGL/Xwx15UcouoJQD5in+9KdG6Dxgl0H8wm9zeYIYayrLSTFrt31KDDdqJupPe
aeW8tL4M0b5/UwBBDcHGkkQUaLWOAgNPmwKhF4y4ZENB5fraRAZ6++rEJIdqkPnu0t+DDgu/K0i1
qFoM38Cv0BhRe8b15q793bmOgLKyGPZYnPFumbbllBKqwmiQzk70Z+8VA3iPtFqf+s5jbvsy4tmO
YNUbktsEXVUlOa1Z0V3Ospl37Wsj+gfbjGNwWc+ESL7UCCYMwy83Xq8EAMRk6uuObnX0bkDHmk9K
OjKZswTlEqT7mfDp963e4Sh8Zbt389f7UGgy0GfkIrvNsawvZ5wzqSMML/MpRPAEh+sQk0pHrC73
CTc+9/syibmh8Qp+r5B9a2IR8oopQwXlqGjw844+LgjHXE/fhq0OxsqXna4QdKRYqlZM2qlg5EKp
QovbAAqz7wqokzd4rlw7ATCtmK18KB2bB+PsfXxu7br2JFZhc9sBQMGX9syauEijRJj+Fl2baSyn
zu/rwL68oPg3iKkFaX73POx1j4+h98C7932hOIz0iXy8Gwnpcn22lmrwBPN/Q8outhxoyxrr/wS1
+tB38lBuSIfRmF1orEbabqbazIogPm0Rc7uO6coWX7sy04xNOkTqeCimZzjAVDjjzwbHLjJIdWJM
b7HgNPKbHiBJxxonDt2Jzj6FJr5BzPEPMH3OXpmuNGlht6bNhC4jy8TX+O2zDSmMLlEfUc4tEsx8
CsEXa4+DBxtNHYWSGvkNPCv/i/RIFBL0TPTdtRux8YcUMk1Lsr4/dYyrSRERO8LpSCOMwP8+o7+0
ggEvqOzJHuJG/qsTenoO9QV9eSTeUbiM6NnVDFBhqIBi6JlJgHZbbinKXM1mMn5kYEAa5oKn8CIo
ykwHGJuBKCxqAVrlnBaZRL05MRbgpIvksgZH6EPfiCX+hhC2hGBf3Xo+rRbB3VDyOenr+ZsLCmv6
+azPgfllHry7Jbx9Th9RxXzEZcvrnNU/yudAcUj0dVkJVT5xGvOA+A7gOj8nvVnlEfKNcEllVuuy
hYUVL9iBoFdeqqjV6Hz0arI/lTln63AEk7sqrZFz10kf8nFHB+zlfqCE5A9FS4RMtz2M+RR0+jkH
bFCIXX0P0ygJJAXIo+mhPLtOKLW/eNmnnkWcvUJRjlewZHVKHPjuadfeSqK8tcrzObHEzgQFmKDF
eTbw2gZtHNrEPBauN1nuxrSjw7eQdgQgI0RtbEYkafLyUdtn0SVFrm/wGJzhCq2m+SzP2zsG8Y93
1EFHqNMu57x0i0wMYgwxfEhoEVjduztzDKNPYSD3nqLbrHvfj0Our5D333+THnOlDcvsD2OE5hr/
TLivixOAzU0TQt/rejM5fC1VxMH6s5BxkvhCf3jMOGR38vwOf1O6gP7/5HTUeYUQKUTJ1wXgipwu
rkuGUqttxFyofu9k4CSK53k9FDNi8ftDMo0X309l++ew5edm/8LjR0DJbP2aYbchbVQQzUdsfZP4
axO0j6TtOnA5yejO8F85Rc4E++eGPN2AuAxypr9qdRDO9rzNmIHguHsfqolYMD+8SXVqZP1bwJIC
UtqSs2rImWWYtG1kXtnLG8lbMy2y8QsIATKvFR2JcdR/bU+wCcrJlN2vcDmrZC1d1BPbFDw0ikDe
z1EOwHR7RRYgiCJG7HDJctxTi+kEiYB4eyRYW6qiZBzj0JO8trknYy2O0mfReuu1dgR9e5ewZjFO
5cbxF7vRwIxvUQ/CQc8JrFZzSLrUsnJB/zLxfBLQICQ4TRHYHvKqO7kPI5CafduBP+kYuXf4ORE4
dSrtPKWFSaE6MiI1Iql/KSjwDiYlfR9BFCFhWFL+UiyVjJ1N+Q5oSit4zSz2YpZsn+a1G028BOuV
M86cGtMET5LhM6SJ0XCsAel1ElLOegWtQomM8C3E5N/8f25uuw+uxZVteZl4TzLm+csmUUyLLkci
p0QiO/T0i5VZEmmwHeHAacON/vZGWRtQMjjPxHD9fOc6S/uLTlKJG6qj6qNSWKqqcKaH5oFwoIXY
KejlfqTEJdP4XxecCA2BQNHrlfxt3LvzskhZj4fX/mZlQ7u5MkNVs/38mYsgSgJuRUHeyJ1YA9xT
s5Bcp2ObCjandCrwzKQLszskfmzgGuLb49Ztwgf10Fdu34VJMrYXjUuUsZBF52fqZPCH+cHZN3vw
+P+GzxKsc083UYig6CQgKHVaxaax36K7G0Vsk8lFRwFKuLzfTf6FcQkGts10jrXu77rh2+S5dI1J
HqCqSaef+eX1vU1LlY9TOVxSLTcY/UmnOeqWminypw8Nbm2TYdJbvXwZH1PZH7tVAVWmLxDomSFx
ORixceeGqWbDA40AmWc+GDx3q3bVoi63KD6rvnQrRrzWDVfQ4jppzn+yYNLQ/p9I3cgX7m+DJg+R
LitOD0IbiROlrDO5D5OJiE5xACcbxfNsxzfFwP4Ai29zJ9ysxy7mI/dJk/rWHxTZhGobw79vFsVN
zfLFVpMWnMAJEK4iUJIVObVB8Tc20mwz9IS+1+VQlxWNVJsBmDznRpQSJyAGIy6qYv+1dNUbWjgj
NlEB176c91DUf9Yu9Fw1QMtkobpZTnVsKlMqjpi3HTUqrSpuC+EQAAeGUk9AT7TzzJykFmWqiMwB
vgyDMFxQ9KPZjQOfhbp1E7arK2znmHE0W19M0QI7Mv2Gkb0aPznGX7Bf65ZZ78L1g1L9JkzQKtdt
p1MQMbqOEWSGAnJ+eSkFTkWohsbWP7uRblkBvYVYXAqGvekieKsvYqgiyRq7bLQ9K3L6xHrhpiCN
0A6wQe37rDeQaTUfHamp7JXXxeU4ZoFx2jZmMUuEyQodWAV8mrSsJpWRQoDYRNT4/mp/9ykU1L2Z
Ah9NG/+QV09U+5RjJpNkSGQJCRE5iY5BhQ0bDqYP9OkINoClH5v9YBFwCAAVeh30qMSeuoIijm6c
O01bn84JjFz+mljK4FHI6g9tSC8/bkfvnlmq99qioG5jE4CD1sF5DH1BgINEWEMrc4IdNDsz3tgS
GHcj9FAvGvvP1uRPvbNae179Ij1qoAWe/LgXUELF92ySE4IHnQtU1R6nMc7++Ah8Og7Pud7Obyhr
cBw7eYnu2pZLttwP9XE5bdeGV4lYT4IhtCYTThQl/K28DWT3rgDVqnbG3hYoDZDiCuFJxx/6Ys3p
5eVff+Izymgwcj7IH6vliboxDTqsKt+8SCWXw5/Z8PnFr1VWnMkaH6N+K0OIdUB5sjXAU87fUrU8
nBAmh3eLjitOORKoAeEfXCFGh5gKcOUKCEwBda3FL7QN93a5AZXV2+e0DerWBqJzMuGTMH1cODNa
OiDI/1oSn8zZQNXvBSuGPlRyjyvS1kpLx7N2d3Ygn+zACJOkLi9zAkIJY1R2IJIXMbM/eyriKc2F
P3kOqwKZWz732CJZ+s7+jwOE5j8qDlc1RXu0he7sE0c5oqTxe8S1Svq++RyKrTAZeTvsLI+Mfn3l
xJk04nNzNMh34U1C4wBZUkoFg9rI2MvPLGRNH+u2/pGBTioz+gWtwxg0JWCvUtYyNWbRpX9Vx5dw
Rj51NgrcRupXHJgQ+3V997fi1K0m3zRKS8ldE+Bqx4WNxylzWvpPsPMoOa06akWjK/Ub3WKDUJy+
6El0gegRVBsKe1ATWsnQenxXGU3HKj9lhBiToGMP8PvuucmzMhhHfJkEylKX/bNBroTv9qlgREpu
nH5xzOts8wI0ugytq9y4R6xtGi98ffrxzGhMnC1SITB41jdCSCGylcfgy6SQMNL+n/B6Xu2S0dUp
+jdRIvQEaHLx1Y5WS1rxipT+vEUaQLU1Rv50mf4HKTAJ2P4aa8vIgvltgkFxbmK4ta8KV8AmflkM
e5jCkv30mJ8zYaJE0xlLD00ejGEyjunBNRMhZgxDbgXoWzzR6avyTrvFSxw3y+wt8tJIEZWaRN/w
4OmN+SXXsHZLC4e2nEARYnWtgBp6FjLA0YeRVwtkI0Thagm+pRhqm0vHeVL+ILD4sBR8FtJyUwtH
hxucXSPhyAoWy8wHB+9D2GCMwli00GbXZLSAI9C3jZS3RX350HeM3FhQvHrijwOoGLu07KSM4K62
GEgy5FHNyGB1IFP23LHZh6Xn/NDBk4CkJPJSO0tCP3OkwlybC9XJfApG8pD7XVwXhMWgpGJ+yQsv
4l6LHhe0SIpKpVyfjtPelofnLTsI0Wq75/I0ytK7S5ZIhwYlFk7kK8pZlgZ/qOhKWUkTo7YkeFLE
NXUGYxrMl/uTWvNaQi1yvpwGc00gHdhS0U8e3vT3LOVAJYFMc6RAk7xIMbEI9+KQa385GU+y2pbs
Gr5YjyKskOra1zWbH7RHY58KCx3cTw2XwD+doOOkZ5Tv24Tb4pAKW9Xrho/M32ey0pcsxCzHHNZ9
aS5Zc9XY4x/vuiYUCuGKg7UcDlIHA9IJ9rQaYM9hHq3wOl1O6yORN57WyQO/1WCo5n0Ro3Kl1Pnc
S994lR8e3iNKgDySPe8lvv+gzW05+a81U8IScgk9huOiszfBiKw/1BVLKLDOBYrf7xr4OivwBrvS
YUxa71+/lCOnIKCGfHDaapnVN4QddAgwAOSf3SjJnnDxsF0rpkW979l3vUtN0oviVX2Ap7XnZ/fM
PEf9BN+0PwEY/d4ZyH3I2ZWlY5jLVTKgAsSE/GSUZXHcsdaydSZEAJ4FDfLxfP5SFUrOgWeY25oU
biO21jvr1lahLDXW8ux11LD/+4ZiIHynNhbk6B96TdC7D22ulXd4XXmZiTgX3wE7rzSdc1h6NA+s
qejHTLdAtdV7BCfKMwAyZuoitDZs1wBdAJawpKRLoLSvQ/M1t0/p3bwqIZQ9jPT1j+FwL3OkPWMA
zHaXX9oB8HxjsbwuDxkHXZuLdbCmTD6JWH54Lm+wERn/Lz1bSiUjfwEhOg6NYJbxI/o/kIynpNBT
0F5YM5buUtylonvZEViDhmCJt/9lL1+sR5+Xf7/nZ/Y7tRDPkHTPHa4PFQ1q2kwyMhc+6MqSmYBZ
Wu6CjH1zMwgOH5+t/ZhYMHNpZXzKOOICtspUWF17NY3nztkQXCKEz/FX8Uk8Ejea9I8p8XZRyCp4
0sBfrTXxjnTyTQ84v6VG1jt6NZyFIT5hOcAwzi2LjkD7gNZ/pLJ3IklTGfV8iT8d6DI9ihVvc4pj
vZ5iRfSp0tAmTG3yHAlpS9LYPEWoJiQoS3ZkVg49lJwx9ORMcuTmDOCSTuAJcl/WQTq8JK6QFE6v
qyTH/N0H+8tjXrKhUkah7+io102u0QZceAfj8AVwSJ5niHADcP+SBUKYgJu9eQybzWc1NDWEuOQE
38csAbfIPxHzgZa0w7GWyWxCy/9vA5F/kWCzKRDXpZwAd7Hi4cdxBoRgrjrfWR5cz1KyimL8keSS
DR6NoOym9DNL2M6VRtYfGRhlm/ZJjYcD77d0ZbTFunx+ICnl8oWYpdE/ZjXcJDici4CPKECSgod6
7hnvnZwezlsag+UntF0dE4OOk4HM03FL5D9AshJh0giqjTFoZ5ZWKmfb76r6nrj53XwABHMtSKnW
Du19B3uFDbDQ1dekwfnYJv/lTHQYIO79GxNPVijb0GAgzVeXjo8N8yNcpccyE08OsKNB0NcZ0sIf
Z0T8Gx4d0jZnHRdzuN6rXf+0fuIQHgfDksfPeQGvW3rv6St+lXm5M364RNV3pXLpk28aAlOohh3W
CzbTfVTJfs0QH3r6KXmD1aBHMu4MZoNmSZVUigGvUoOzJKFfh86pb+i6v+Dmc/ciVcD1iBnva55d
GSvFC82x2nZ3MprEGi9YOKiJ3AUIW1lh+XiUWmqQjhpnoRhpNikx11A9xiC7dwELV2z47Zh4vZAU
GaKvrvWrg7HmWxld8hRGbj65QbaYUsP+TZh0GaSwR8Db0h5x8ej9El5PGlhufEWf9LeE1iQwzdXc
mFKCWy6FlsXIS/JutXDaHO+WulWVcF2MO93V8Fo/JoxAoP0XtVTzlK6IEXxScf+V4Ru4e5C2x5ZG
/9kF5UTxqNOrLVVyPBArQnvzDOwW91xBffARPPqEm85WjBeaLFLclJ9zqAf1AfSupzXPQqpLl9c/
LcEjaCCTtYhUqPHJkSgFJ+Gt433VTXeN+mOX93tgB+tRiObfXpcegjdjsRmJ5aORqI9SWego075z
ZyLh9+W0H8luiWg1v31zpV/A8bixSF90a3Tz6u9hbgUL0scnsDpWdxCrs6/Cz6RTNr3G20uCj2iN
HDc8hfL9HzS/Li0wN7UI3WG1fOQYooavRFERVcFXwYYSWwLqWFnzPSHR98//bR5H2KWPPoG301dz
Ku53o9L26u4CHnsSraiwPWSqsJfX3UCubEhk6pLg0o1Z8pshPZ9qMEbOOMzxwHe6ItET4XNLsfGZ
dzAmIWE61TgPiXBAQIEP97dBxVJ7QrkOkvypkn/EBeaVLCzVdPJbGpZpPJXPgZhgV3upz4ldl2jj
FBpuF22sfMB8F+aUwZXKBft3w4QAhLqKI+NAU0Lms6t6mq0V9GyGLlxjQPXOOtpE0XSywsK9mheB
UGQE3HoYGukivTI2jLDibN+h9y2VFOAlsbGEEr5J7ILokOH0M2MI1oe+LF9wg+aCpUF0QwAMFYVw
uN8geq/OWAO+RbVhmcRCHM98NZFx8FaFWtMvBEJS2BuL5M326gIQYgZb9WKMJ54h60YDmaY7PaFs
VIQq2sbNdD4KN1bfe3T45TRC8wMWXigVnz4bXY7g+2Icixs+6zIC/4CGxYuEAy5zVaxPh7u54c3I
MYJ38gayD4N/fBn+rb1gtM6pAWtgtqi6qlESCXW03aEBDy/aKZF082fbHTeM0aEaxfLiSNY2pe+3
zjsUIuhkgRgtDh1KZ4B0j2u8U24pBfOHSCk0uZfvMLi/dFUeVSNe8VDwlFR3Tm14mPXbX1gdYFn1
o4eRiz3zMyNuUHsbyZSzJMNw6R1dQymj/V//gvfpHtUwjV9lHmPyR3GMypuQeNJXMCdJJC8srZvM
FNBBiLw8YFp6EiwgacqiBiqqPNwew3r6NXRgVJwmYphUsl5BZeoQbWS6I6FezUeOBIhJovAyDx9g
yPbpYvIgMOKZ9ZoR+F/l9WeoMisWDuxew7saizZmPCmcG25seLOieEIJaeSllaVnbJCLlZsE91Rb
3boyt+fUVBc/ZByCc3QbnjKfbkXtkYnEpJKBZBAvWAmPGT1Vspv1AMwcdb2nOatt/Hm+qpCol7vM
3uB+8VgeHQUYCKvv3MNltRdbDzBNLdkYg7W1ABy1NJKXyGw2PeHRLOAXgSFIqE4QPFdiN72RxZpr
Pv+sgcKf0rX/SB03vyavdk58nt8XwoazcPBeZL1V1IfNGdUlPwpJn7p6qe3WtncFGlh0uh6DSIfw
uJMDNErPhj2woJ473HZA2JfdJZhmGQnv3+AEq5hmuZgasIDZVH5fITTCAwd4XP2TO7GLB6nyHK5Y
8Uv9IlLZdpDpUwMxiMJUYwlCA2M+W+v22dMiEkpzlkt0r8/8PUhNeKgx9G3HREuPjXMT8Q+lryxw
wJnPYKdz1LCF5IGEJf6BvrtCrmWAA/lBeaubcDu2fLIj6V7dJW0VK7w07LLtlbMGNMT3hiQ6LqzF
PTiL9EhoXuyHhhxgqRApAOvuQwzjgKX8VGw8meLzu6YCkcWphPZoxC4DxTdtSVlJ8uwxgm9gprwo
+SaYcwqJhl4WcPyxezHle8iq25atAtXXcalu58sEKiz+YjsQEQyoDtsXtuh7mulF4Y84s9HPXWLF
RFRqt0VHySOMRmp8Mx5JRlvh/2WGxMfb+HcpDlG23lsc3lCKVVkhNXwWAx0FTEjA65R63hRJLkUg
TDxpUagtA/N5naoMZY3N7FZjEewayIGiP47TWRxoINu6W+g67+vwjjfEymVk4mwzQCSk7jQIZRoy
Hj48k6PEl0aL/BC3XLcfIcj5RFFMKtYbWwQD8PhGWGKAx1xrWhIIKWSdt427NKdalWnwXsXco8Rm
D8/6Uv4C3k+8VztXWD+aGDoX2EnogTjljcjhX8Bfq3TPwm6CRjh4BB8qlz38wDi+XOE+DeJYkyhG
IgrvsSuXoEFntX5L+Ofp9jg0A8GIS7gRkihGeWfNH3xQqCH2+FDSOf1qScIQygHu2KSr3W+PB2EF
D98qO4oTqXlUJULpJHjFRvYmh2uagdOgw39sVe0zOKybwOrokGYFWbTJUWQ+r9TkqYgjLa8bVZc4
+zRq3kEE5gGm5SVUsLTGt1hpR/Dmv4qfGjC0+s33IaZCDt0GPtFqnQLPZWmy42Fcj8fNux9ruozJ
NWGFpAbhU0w3DFRhQxz8/l+gxUsxsLfQhML0AC4SaMHatRtD16Eq5S14Rf2k4kFfMBmbbQcEERW4
0pERcVBjHmiAeP5zwT5hxfcbO2AHR2gjEmSF1Sim11qtFV/WhN7FrCOW/hNSTQjVQD25C/qUu/Zx
aCQhcZyOtTLhY2IK1n4hrZlyxY5Ofsru3Gkeq7re7VbSmM/EDxYHSGyVHvlhd6gHcQXJgzMEDLNk
kdZEdpvosubEBuxk+OcEuBbchVy4GTezQpn8zUePxj/1GaeaTrTNjuu/i6JOTnho3YG4gN7FOhCw
Xt4WpPjpyBarsX1EBrXObvFBBtOGR9XuNWgf6GArgqeLaqPHoJKqQERzAccEkBz9NwGBqCAEz/Fh
Dn9ndebrDXsY7kQ7bLICo7z5wrWMZEN2SvSNOAGWN9N1ExkYH9RDKpRQ8UG57tIAvglHNln42wFB
/3NTl6jostN+24Rh7crAg99h2ixDjzL0Z9LX0Bv/Now8sJzPmQioMgXuk/Kz329gsz/WmOe37/BL
K3M0PgcEwJhdzfhgTaSn4LcLOR/6ChI552pyLjeVSwYlBgqKSgut/p1vyntsTtSlSTfeqt8liACe
G5SRYiS5lpQ9OlgYCDCQOuotwTaw9KoGxlh32aKeLV45YsxsY0yuTBz6gHGH9EXRpXYk6MwIC6TD
Td76TEPmDnHpecdn27Ld/3h+4nvRFoRjz3+DeqhQNjyGAE9zsWMOdNWCDrG4cwM6vp4GGv3ejZGI
9P6mM4S8zDMCbUxidHcPj6B2XJxPbIH86rUl57eatR/uq83HNbrilwuUrWYEUxL9loCqgkFko6+D
zwA9AmFu+XvEU0TB+3HDUZ8neKJCQE4E5N9fwYJWc/e35o8YIxVA2X5o3Dj1SHLTRVuT2e27JEVr
yv9UpsS0IXmneLE75dQSuhTW1P/ASNintqsXxnheFIa7Cgd1WfutQlW5HrRvPED2vVlv06zAgex+
3MZrnJ7Fll47p3nHwQD0hgGHip9S2IWM47rhF8LbAbioLYI9Tz13pTf4N8xbWrYA3gL8UnGuuFDZ
blMc1jNy0qHxi+DPJg/yLhFtCry62WRkde5XRfodRGR++vsyIg2uY/lBkA1jjckTQBuHX76Rt4ba
0oxkwUIxaSdKaYsVZ3E4G80XgeGXb3Yg1NF56Oa6LnFMZ/tEWDv/HFE5WSpMGysT54/4/bpEYINl
tt7BV9byVABz6KRWE4a98fmUDUhUFCdi9XQkLTV+AOd8QR8d/OhrzapUnivhq40mgV1MRsr5NOW0
11XNxTbeJ4jauc+/D6Zw39BQqSUjnulsrQxexzP/TUoKsjAGzI3ucq2cVcFQfu8WpPT205jfAUlN
O5/hfsKos8qZ56KXLUk+r7hAql2UAi4q//wqtDI+Y+LYgvOfC3KtZKWlTe1BCuBfoljG7slaXMJG
V8fEJeq5eze+irpGGDcGZ66n6URwe2uf/jS2ymgHYLXL9pcEqX2pq86UFBUaetnk/yjTfHfAHX2K
vZpeg5wjX2gzcgQubAgk1T7V8amBosKEZEs1b3XCDhmF5vKF5/TyBdRFoIzg2ViToiN2dr+kN7M/
p/o0sSticp5AuaS+reF2avp5G3kqbiTkhkc2xVY8BVGlhe3o3KWhjwAZZktXeDbvbW8VNBl8KCJH
9TAtz82Z8+muRy5CgY0I8M/2k7mlMpPmiysUAAiaGnlWivp+M8LaWoqp6NwiJPqE+pXzeOwolll9
tOT/91tKMnM9mcXM8S2PnJdJnBlZZJ91qZTCBwi18cn0CsIIIwREDOxYTqfzhWdhnbMuVE6Ch8BV
3sLV9D7GE3T/gvRjI5XgCSzO21bTpSO8rWt2e3+a11rSc4LXDCHbn4/enQFPx6F6BFN7y3oTimDE
VWd63UnZikl1/uMYRK73n6/VxmWrmwKFttfvZA6jePjJwlb2mm/VR7gW4Lpvjf/qpdTqcYv8jxic
MSOy4asNv00gBadnqgoBwzjdSuu4+OWaNNvrXXVIdnBIkkMUxtamwnDCx2IjSjIMuXjZEQ6JJr3B
MtAO7KSv4E/oBVa2rXxnWXaHc9vnhkh4tnMLXH9C01F24aMEeVa5jZHRNPHqtuxPwNL9NmGLKTrc
zaUEAMC63kyRz+61Rc6eUY/nvSDmPwJWfpMX9zDNNCXpm9ZLbvFhQzcy2iMjUq1G+hntroCFycdr
/3mvxkb6BE4OVYtLFnIWXmLBrpZX+sCZy1vX0F26XEV4+IRid3wz/pcokvl0fZesxyduX2OU40R7
oUtYwvvlYv2DtWqA1stUM8gXDZFON8cPShl1eI9XetpqOZcpBEtEEpyd3ziNS8O8mIk2AcbivoXe
3bSzm/les4oY4/Jkwftp7YJ5TKOhfzDsSI1ATQH2GgedU+uj5Afzez1/kvcwJGK6DaYq5o5Y0wyQ
1yYlIkzjBAuyYnyVQxik+AiKDI2daSllkNMKDYuz3mMntxCEy35kxIv5x28Mfnt3THMiO0q907Ki
uFqYdhGMFtOYjtAdnYlCHuFtALCQA/hEg+LTZVGdfBz4aTPMZFbfJfjekUhoRPWVVCVjBy3JfFrx
gfKlhIsH9fJoRIBn3cyYtLIcl3SCq2fhaiwy+zI+RlgNdjQ62jQGZDyK0Vcc27u8Ofy3PGuRPj1B
hjc0/VDy6lOFlNo8nZHgoiCqgxxuwy067i5Bn9Z915g80lHFzxnalp1MIeVeoDQBo4gj4wYIP9Nn
yqlziAYZefCr8kjEQN7dUrgDF8lDN6h69GM/elMCQuWDs8stiurpmTL+105KroH3fRuqLjWMYW9F
BnV0xFSAMOUL3yOGHkuyrASxg0Qx01Lidd1KzJdS/KtNxR7AqG8m15+UWONJTzcsSuag5yo4aahj
Bp/1CFpnSGwIZOv4jsQFI6ppEnirYtp/olawwbiPjgjBQDKHrQZyKqzE/YHeganGJ8CMRGSHE5vu
Mcq/dXPgfiMbqrlshJjmNd51VW8JaSKKUsz7Vtpc6/IMyEAqg6wrkimdtMJrH0ETSfWNdyBZsxaQ
KJdc+O2gzzBZvpcg6oiKkHNrDc8qDZbgn61MAuQ7qbs+byJgUpXq2pwa32VPsAyCjfBPcWyNNh4w
XDyS6GVLUNfJpRKSJB/a5ZDSdIUApOeUIJmWVT+8q3iodW6GblgKSw9dimO1C0JSR3K26impLLTR
jnL2TGMQk/dr28n9N07nmn5M+BVlKBRnpNclCrLhanXRTciENwd9raiDa4l46gksh9AsmD1TFMJY
1aAcvT3qkxXkNj5V/rdxG1ef89GihiGbV6zCEa11LzQUV4zsZNUUSvWfm+My40XIQ+FXNEggLkPf
ftw1EYvaKU/P7ZYrpbTh/fHla3BGcbxS7Tto7o/67Q6/xcXcv9qIIB2nsELNdZYx54Li7Y5Dhrk9
rR3CaoqjQVlagwXuxvFDoG0sAFktRSQgce9fk4uH0k/mTE+xNQPHbii5Zf8YVkXHEEEwKrIzaQ+g
OFzsZUIhCToxf+RAok9qadr/MQtC1wnPKww6blZ91AymQEPFfUHqVU74OkK5zGfdEmBQ04MOnqFe
COJNPlrlpYKMIMV/hDhFVkRlG2nnSqvWeJe1JdswdCcoxZAUn+vPM/DEGhqBf/tt2WkoYfm2Yi+8
sUAnnVf8KaYkS/XzpeK4aoNys3uwIopAtePXw7rUx+glD0UpBsUYOja0W1YQU8fBSzLQVkTWT0Po
m7zZssaG04P7jN6OpgkOXZJSGhrm9oJJLD6Wjy7ljHDECkaF38KQfAiO9HyONnOYKEEwRC6gSfXu
HqoVbLiBiHr88YqEfNxJPR9rLA2ebtVx8YYuI8oJP+/pq/Q+Rp/SkJasgijxAs0iOquX9L6LC1IU
PffH3yrzN1IXZJu+/RlIZnIRR/boYH1cl8jpVi1XuTJjsN2ypUgJUuqTjUoJBKkfmIX0tvkpT6HJ
wHfsThVWFB8j9chQ3EvPTtoWSlYQfFNxYchbvYBGJUJY/xD7tlqLKQydsRlgygjHlIAbYCf1D300
fDUQ4S7JTxS30OtvVhxmAwcKH8rCUX61RyT03ROcLTqRMDmlDXGw03o65fCyieYrbmnJApR16+QN
+SIXsXSs6spt1twpbf5hTXAcxEtEfeHNPhw9wkpXzCWSRZ6liBHDG8MNOeMJVCU7lKNzY1k/3ihU
MLbHYI651WkQce2G8C0dGTRsU1doWjLKSX6cSEgekR5Kh4SaRfDPmoVb1RYZESuIOO8Wr92m2tL9
N8EQoLnQ0KLTOAaUMdFxLb+y0aPDfDNF4uGnePq7ueyA6MbmDYwIUmoRwqBNvBGjewKCkz7PZM+Z
UM1ipR27VXaDe2V6n32kMu0jMJXlPth0WSFMc4v/iqiyNctrLoGImkMKQreAG+EKIj3NBsw+t/6I
HUL3hdDbc3SP/mAq5PHJX7yTh2JnrnncgayD1GHTEMSL6Id3XgtOMpuyBhNKv5J5QCDVvdmLRstu
veQLsLnf5lL1faMTGYOYiF/YXUYZse3rax+S3UM7L4U+2LsHzWUAYUSsVvB/IIn+7MfDP+EGO5Sb
GKN8KsBsmBYHOpOl+OM/Xls9NhJQFe+hiYPDErdaWAssPUwq08bqfgGDAW7rrjrcG2lzy3gzfzZR
GvxjS22RA5I5hUx5I4+fXk/Do3lvFYJ4IwVxFFpmsGk37/WEfAmF5WU4JOJ//8u8u2eOjC+OYg5H
1pvWPZXcDaM1kTU5LCB+B3R7TiFCU6SNyZgHH/jojx+m/0BdsK4C+LgRaMPy65iTRLmx7UzWcKeT
1lqZpmbHfOOOM/4FSZ6wa7NGvsFhghMo1UVWOy7X1jsod2FTmJJiDWO7NjK68yM9Zw47wuNnmde3
X59IRH9GvE5yOobSqOKX0DseGVzd6IMjcWeDij0G8XUUhDuSayJ6Ifh1KZLx2aJOiowAVBHlN9l8
Cu2o9Ji2yctbOn6YTC4Pp+NJ7E9zgvSqRZbA8cds3JxbXc86YkpIS7QAEkSv4uf4wGjPSaW/+GGV
RhFEx6dmm2WkzToGIypeltVaF8Ja5YRIwdknRBJnP5orDv+rW1B9sjAEqkfGAahaIsN2QkVgD8z/
+L+58zTfz4pYbfMlzJx8DHGmGh6V8/PFrYojpsJuqCoMzSyud31n5eCHLVIFK8oIBecmZeAFW1QU
e5QW2UX8uDAkVCzOh1ZBJY7YkIf5yK6uWLBuaDE77mzMYa/hS4lLGaD3szZgZJDlP92BGLvjWfix
EwXgYS0A2vKb11ssc6NAerMoVaJO+Z+mtKVffebbK4D9DEODHM6gROy60uVhPNfnD1YMHVLG4wy8
tSSx0x/wAB2uZFUD9aXJgGuhD/dzta/lkTJ+oU8u/M9YUGAsKHslYAhQvILUwZA3Lu31Sz3wysVo
TrCT+QmT3YMaZvSEeQMFWiCM0DDjsHZsFHTykT76Ma9Dvec4+5B+LCgq4fpp9tJhN+hcJCZ7xeDy
AbhjGshHac8R/m30EgIqtzO6k+xPLjGbC1TrRQlw4gzfDBvVY3CEAzxnaG2VvfRf9KjOoVJb8HTS
NO8K2VszWAXNr980c70bG3nZ89prZOQ0QRCfgcP2oMew0cmhuauqMWL8t7ErGrhcXTIpnUSr6pmp
l1IbhhMl56r8hGFKksblrmAwzKXTk9jqnkbkDq3j0xT65nuYGX2BZeiajowlctOAuWCi2fsruFve
nv4Dr65BvW2mGNCzpCAK4rzGIq0DiAAkAyRsbFWc/BZPP+utW7BdMtAIjiXwDX2v8vzrC9aaQEH8
ERF23TtdMF9MOjcJli4hOp8ovz6WoaNahso2bf8rJjuS93zAh4vEpb9ly1bmDmAVxTUdq1ib7rZw
PUQBy+slrgJCuVQVw3O8bSe1iX5H4XyNt2w4ncQvDXG4RC66Egar349CIA31Dq1UmmpUaEYMh9X+
q9o1YdQpF2oAXggqMHfa/0W6AMyyHlcFh+W1r+rTp1rkn5UgabnrM/XVe+66y9vRz/0hsm3tI43l
YX/+jcJk7w3O/mXR1V3+ARFp/YPbq9vtkC/iWV2XcdCQAJvzV0iR+bll6qVaB6vubTnbDZ7n9COK
jjmkBykGotZca25K5o/k38dTIKzc6x8LRYP4WZVM33F0LLjibX8xfW48EOJkLmXQE2eT8f20nmUq
l3vYOFIB5gFS1m4ptkcRUhqnYCEHU7EwbMDpw6vJzGEcpqjxltUTWIcA1Ce2Ee/m0Aprl80T+y2e
k6pz5QQQ0RXIJOW2fmAGIYHswODmRxoaYOuXqTPqOcePr1aZS5dvR9M2kSgupej9Hu5sHSHV9Ach
0xYBLz/dE47FZPKKeIfB9TtyDLrT244nqCWen/aPQJqIXjsr9EMYpHu7g01y8fu5itnia/FRAY0f
fr+xqUryf9VRmetpDgRaK3ao5zbSPbQBOhJMyrlf7zTvv6Gu65gfj6w13t+W9KfP7tERZyzZXFGC
lhbSxxPRdlVwyN5Jo9xFWBjxl8wSmGU5Ci17OLlroyIJFHNfRjEt34se4UvsHawJEVUi5pja9UwC
mo6Y8YtEtiMGoMN9/BLcceHjgQ0LBxGBdry2c5X73uDgor6RG6IFxw9EyO0z3A+h0NY7UGoX9jdL
wCaXT7chNRib3IIQsvicEeOIJzm16oLypy0jFGU1adVPbCCAFw7H0MRBewgiuKqy5DyCPuA/dlLt
9/2wtETjTaIRMYRVRXu4DH/pgdE7Lp9cshlDiDKV5qkE+DYa1a7oe0yDLInI163z4dRZtp2x0pgq
ijMkuITB03Ur3DaIIpbJzneCwoj5v5cb0CwjVne9LnR4KKn5NRf5in1LVAu5pHQrT7Cw3Bf5tHT3
JERZohnYyPDKJfgYvRMNGUxV6LJa4K7ceG+owhRynxaPE93JAEiIeUEP/7KxH0wUHOZ6xork5eAc
bXCoeDfBb8ORNpRhlqu38FzbtkT18Gj/hurljW5b4u6JeIadBYaC3yKUj3BBO31f0KklDN0SXh9V
o9e19YitowvjodZOJ9qeJ6C/ztp8IOj4O0/IVS44vR5X89DG0HrFxI4xgBWw5NA1VXzWF6vgvJ6G
ITgDavgw6Miyx/aKgylbANNPHcf4kisy2zT3Lm13kLjxIkGRcivSiUyFhdPwafh6us01UGnp4E7y
HDxvP0Q1tGYwhbbcfpGaCnH3epBYpx4Jc7VtNqVtUK+psmsF1lkmg6BIemGSxVtV6/Psr6egoEoK
EMGYf7mD+E8oz63IMzJJlqMCGcuxSZhPNUSWQxs7+xD/2nQMj0RkZLuxjHUhLNdwrg/8WODOiHgv
UtCjNP08Zskw7o3PxLL2Fk6tijni6yE859Z/HnTb4R4PSDlFxNimH5RUi3YQPMTZnbOdhavXPDGI
k7STwLTPuHy4m9fUlHIM4RLmdhP3Kuog4zbyZabhZFX9c2/Mlgqv/9EgFTw97xtWRaLtzXSed3Bk
b5f8hhIaTXLg7SZTl38tK+iv3gKERtxNvIwzo6IF1oTgn+hO7EsGB65ZlCweFcBIGVK3mLG0nA7/
PpiDHOgIee1VYaxzsre73jLln4umQxj9HubiBU5nktcNoLIzpb6WE1VNuvr6ro2mxSgp9XbVcq4s
hSjao9ooh2IeN/69xk8UijTfyJXiJPiX1ZLVVH+eX6m5zVvQC8rxP5msYz8TNY8KCVslx9GWUF5O
70Nw13uJB35pApxWKOdCm1bgr06vBPJ7nG2/LnB0Z74hFOjJlMPK/QcRwKet80Y/DlfevGUSrVU1
9vaKaMTTM9adEI2U5Aa9FSEbfhepJ3UqVvfm5TLvRu/w1rmR0k83w27IlNVX+kOeZJ5zUE4HPgh+
RjpjfX8QgRvEHRdIb79R7LWZK9rvt2g/3DBBJaAUN8v/2yS2GnQAKYlKbVAlPunTe5/RZRU3+8ad
Wmx49FQrL+/IbabhFuGVHVtBS+utB3EeiZsBMwoaLuXv1ttR+cobqkZHEAu8qN90J+haSlEzTgTc
E9KgVup/AtycKfpE2AmYaObAcTwNO56+iPCZNfJK3IlBch9xDUMtwaV6oMLTayN1Dn48kNwPvQoG
6yXj2JhTrKG4WsBCiMsw5o734z29YW/lMAJuzJViMzBBrlOFPcEVfQdTxxD6JkxM575sPeKusUEl
fXPmY5aQsgEJwWW1cilZDTumIfVSe/EW0d5+xNlvAxYuA9phJ4Mo+255MJGg/cJa4gpko0quzqMp
ujP8MTUPWySwkjxOZL+tFlshJkU86trnpVAlWlLEvoISOF1FQ7DKQV0z13IOVVH4tp6RAs85oEV2
ZwixALinyKrgGUKSk0NGT9zVAucPISUK1yLoEgmkKWj2zeTeyr60hRV62JOivHFthyobEpV3/vc6
QeTePY4O7r4GacS7nJzzphvm8K97tNhoMUhtvXWdXyqkgXeefl4ZJAN5AcjUiFGpb48LFzDSKedJ
kOubq/m/UzafcC8yHpXnHOlB578A+6nPqxEZgSHrXqFIOopf5a0Q+2R3u9tv2mf7eM4g92LftdoO
7PwkY1VhiFT3gIu7Ftz7GrdQrnc6obpBHvqMqOY8f54ocgve1nKV710QnW6g1428HHPU4Av1J3SU
aEAw/u/Pi5OQRyZgGpxgF84jrBTgKLG2j7wjTi3j1bdaJoP2VKuqUrcoUb8mTm1tBMFKkQxo7SR5
mx9mFtgy45XD7CEjBl1btZ2eVGBMSNGWlMEeCfl4QuyP3Lq5K17pwowZs27HUn5Y199u4ph3N7Jj
KeXe+OW3l2qsgD4QAYd19SmGFZDHTxKDeD9rapSLosUb3vVUSefI0ueyuprydCp7cy1n9ck0re4H
IdKwsuJgR7GrPxwARNbMVkRIiqjo2f8Fia83URZRMmwSzszqpIS66azYsurZeBKyiAPD/XFRKgAS
0YpaZeU35xuUs11L+Bdr7JAdHs+QVyG/+qbmbgyW2fGaiKPKVKzwose+sQhMGHwxIWL6pZWJZx7m
oBFMNoxVKQvMdcKnRgb+W8a59HyjwNjFu8W1QKGbG8aCkQWXiNk6em81BV8XDr2i4yF0XWosKqSk
uoTqkSPxltdAOO6yEQF7kKJtrTUewsDNdYzFwfgMoTOPyUCO0DXCtQtUKpJ4ky2QejCpHQ9Wn7XJ
sgQcow9BoPet9h5EAs+vdEu7B3xuQPf/5IlIw5V4dOhkRoHgnGM8Jq3hVpWksFlOu6IChh9c3jx5
xkff0A45jOKUM0Zv4Hq2FghNV0zg6mvqaUNs0U9FWzFOO5bZYFQh9ale2VwFtCGdZAk69JIsjfqv
FtNjMCvbntwv1sxcYRn8y5nIv/N7sgbL/YqBf0BgkPRWo34dg+GnthYRX+Duh6Lx58flhT0eI9SV
Q7sq2Ht8lJvuSq8B64Vc1vX2Y10aZiKpHXePf6VfKdx3lio3Ti9k3NIgKU5zA4pNGkOCcQWQHIuJ
kXQehA562ziP+7F0s1W2JISRhqT6PLCJo71F7Zgn4kXKhhNk5t1RFmePgaAhgPcdtIGDEm7LuFvc
7g+lIl8Hcy/GEKwSPAFt3PnMlY17OJr1416ZWT9msNoaXdJaLls6SLvhwqJmtxtScBKXkX0L7cG5
BYMTtdARZ3+ZQb1F5OI88XG4Fe/HWBUGc85juUA8Goh/KjnIJgchc88oEj1TDWy/5BM8+Lrv1xSj
TuDgxEMqmq9nRX0i7wHhuJYI+MC0F0l1PdVKIgK4aL/VoLpwT6vzECR6vpdSrTM37+86wR6gcAMo
7BJK6NtoAbQYresHP/pfwWXhjQs3xzhy53Gou7iHxC4FMDdmwcDz16PuntfuGN/VZUfhxxQPS6se
rRp4fCQE0cDCe8YePJYsd+5bECrPG9XJ0T87nZ12K53B8pGVYI5Eotzwba9sZ2fzgytLIerKQasc
Jje2CSA2wr2v2SFuUWDjCRoRaGqHMsB3U3TqwFEUxu9QLx7U47Zp8Nusmw8BgTMj2FZDum8CTqT+
DcFsKYOwSHjh61R2BsLILCiQphjAE+PNV5LN8yvDp8L+Uw6FxHXkwfFtUwuWOkPeYt20qhqwc44D
/pVuY8Iuw2H4y466itfqFkz5OVFZm7KqcjQjgMfI3HlZ/CCcBo1Kcu9dz5vHnsD2v0BclZsWfuuq
SY/dPDok+7SN6AqOL/cjO5fg768P4DvWYqz2zWmaTWSLJq7tulteapss/cSS69iaoQiC7HBqwHRZ
ki/Gmez9qF9HS4613F6y62Mod3ggMHwuc/OzJ0uFz6kax5L29CpHoK5IwLB2RcTRi25NfShALqdv
BF24vjiIaEG+j2SJsptv6MypOjEQxwDa5YKj05JjB73YgO+wwBAsu5JKAB/KKjfuTmnDkn87h2ZD
87O8Uhiuavvv2dL+fKhlBgnAp3beJHzvSXvMyZ4PMja3M4oBiuNhes5HTH81tuugOrGUfsO3WvX5
hupUblYXoPJbQtt9loeazNRsuDpudpq5I8WotkSA6XeTCPnOGyFHROvvd7mlxg4wZQQJY2178ng4
jKUL5TsY6SGa+wzyBI4MfGiPHwlhhNmL+VgrPy3NwAaIgqecCMBJD7iiawrh5UMdBBftyUDH7QKf
+ovImrFbm1dtjbyoDQqEabZ69aQEISPBRi8w49Xwis8DnBJ1dA7gdwsicSsazfVpdw4w0WevOHe+
IyXEx02dN09Phuz7PuApJ2qGrnTnDopyG1IPpJ6kreSMlETP+pzCaQU6wtkAHyVrABm3K33G+9ue
04KOmghqAsdEhessy6WPeKlRfPweqxq4PF+dCHMWXUwdLiPgJgvlCQrYquhXEXzYCsG/NclfR2Ra
iGQvYHAFGvTFvAXby36RwCnFfMCoK2uL/M28j+AAvHclpv6PsRQCg59HwphciCpJ+3BYhAbnoFsk
zUeXtIqFGCur0a59pQljyexkXbXDUmihDBZhErtfs2Omtem7oXLTt+bHkaacqbfaFkXZu5s39AuY
lqEu7uyDZA/KCSrYfje4HlqqR5ViDkvb25+9k45qBECsMbzcjlfI92IkXta7dxVFTG70hlKDK7lo
5nO/5BKAscQoaRtd7uDMxyeSL5q7oCYz/4Mr2NYmrILmroIOTmfqwihXYU6S0yJDaARQRaxeOEhD
rXgumzCYDnAXUufI4nGgDtvaG1H/mbKoqDuy2DUiOEXnEt0NRR99UNzZ9tE8jCYqWx6elVSaw4Ki
Q0442PD/sBTNCsL/1K4GEzUnq5Eu6yvCPjb0YetLUmvbAysl5N2OQOfmMCb/ntPx3/gqdpW8c3Gh
W3l/brA42j2sdl55+Orm19D7nX2oaz/wFFKOhcIVz5kzOMTqd++i4EyR58nI/3QcB4/C9AOfXPnw
yX4j/G+rRHoQUJBRhr/GFpNZ1W1fLjEfu7e5ox8cP4Z0fUty8zhE9TBsrwdfBV46v7R/UlmViVhN
dodDEzUjqSaNwT7bpjG+3Jr2TRrmrsJao/5Ofdh8b8tkKHHUlLmbuROVvO1ifLrDH9hFb6FUHioe
wm8VOIo3pLMJiaJzIlpJRcFagIpGK/JQAVWpFqVFgE48FLTbRSLOtpu7Yl3njg1O/YfUm69sfK7A
CIlNx2sgxCltolzUeBHNe+rl0TNreX6+IQNm0kBCA+8Cjh0YFzc8ujGBEHZ3PH76S9u7i8hRyIxw
vUyorxtDDA9/lhRI98ow+IkG1QnvlWRTpVPbX7kMD2JU46SQ2xLztXX7DYQjw5eyBR8/znuFTgRW
qCSJEiKVaReuUrJe5DjnB5eLKg6AF4w4qS+sCN2dGJdlrk8bg3IRsQVMQHOUa+/lE55UXbtAGozQ
u7TuWMCjOcULeNikuZzcJEwmAm1mH9fZHq3e0yE0NVC9xtYd8tHBL/jwMo4NHwk+8pn8PKOcn8e/
RYf2dckPmghcafHHk8wQ1supeWkSrH6Fx4YPnJkbpBieDt0uXBMe3N7sQpIp2x0U+bqQMQcj2+zD
UqMRbSXIAL1r9sed5qORNXnbltu7n10vtyDLugWiVSkEMhx+QhWnKXD3rPovd8Q7GhTQMujxT/wA
XolDQvUzZZjwxu6y2PtSL+EVMxcEJnWLqEGtr5U0fsu+tcac0X5pPvHCb0n7ciWb8gVDf1PrWnLT
CV3M/nTw1I9LT1XZ2KF0Y36L4seAZpEQoYm7Ul9hVfVCUt9O8X14Vqm0OozMkNu/33WLSqirj8Jf
h/w2WUP8fHrR+YT0U1qBoW1FB18EAtF+kvnbnFcZZ71ez5sISSj55myJ/TEYvIwdSMpB0Mzcd2d0
FY3q3IlxNDxjlytcVGmZi4XLh5y/Oey8DgI0FTMFkALehQQEwKW15KDp29kntV6lKcGH406kYsbx
P25N6vQUmVwMAUqgZw3AfSdhS5GUF8R9M+vHazvToe8/0d5BBrkthcEeBCrhEDcw0eF4aRLkIkR7
LHYgv3vmdgUIvIRRTz3FNJlbR6OZI7cMAViawBAsCmq/SgfMJiEd2gATad9d3M/sXfVYM+8pT4LY
PnftQqm1XHpvX0LHbqzzE+8BMna+3K+1mEZGk50vNXuOhnWETG4KQ6OTJUV0z98GZiaD9tTXAyKp
wL8PaUGAYh4tdRH424OyQInWeJgTIVGrSAVStYeNmw0bmG7M5vunLNmsagVkLr08OAMbSHardyrr
4BlDGEdbZr8fwNAWDJNddPyIMhP0lmFDtfkpGYOqdj9iuDbyQyw8PfOJEGc8AfSgfZjvt6sJRA4/
10JkJY5lCFAXY1fhDKrLYsKP4jUGCqCL7WIX/6qeXX+yMnK44I6SAQMofDZd8Q/drzaKCJcS9G2P
hnsTpH9M5a/XCLVdwPUtGPXVJ8bRDO1XHxbjXAob+5OTL1p+YfR76cUFshZiMRqjS5FZdt3dkbIt
0t0JrpZkAsrLFPLS/6lRzhusdNvV49ZoawJ+Hxo6fgulUcRizShsvA2tEN2Gz7geEaUpf/Opdd/p
29Vwt/PsxmcUZiT6kjwEgtD662Od5rR+f5a1grDKNKEO1s+IqdOQOrrGbmgxznJaIxrHDNoYLGaN
bTnAmS8jpG1qNHo6VGN434YtBXLryNpEtQWONFg21G1R1iYyo7rKuX71/x6NSGrcjNmk9b694MYD
VDy41aAboLuQb4IY17Vg+4a2MPDoD4LdeXsIMH/8XRiZ+uxDluOJdG0YuQ/LaWhecdEwnue0rEpD
hMPaNxhX98XMXK6eN5VhfAc7gMR+hvntXhWVNQICcLok6S49ZO/mQFMVvm22W4PPZrzLbpGOAhJ+
OC9ytKuur4yIQadML84ADCEJJxKRP3zt+y4V+AWwHjK0D2uTnBqRhiRMW+owzixMkiWxIZyjiWGl
cJG5IKcrSFdDgmPgXLwPIbmgzuYGKW1kfTm8ssavc/mU4qadMM4LArrKMWD4KaR+fewM3s6ld+fp
G8QYMxszMfrdaBcb4J+8rucm/W6/f+phzW8uiS7SCcAs/58xoUlNylYgXibs7Ess4OW+/UlKuGCh
LkVX8b2h5Lb9JCryOtM2FVAtEJiYfqo9Ga5OPUKGUtfnlrnqtvbOyidTI3E5iYFydofZGdfr6ECh
kKGqokxrOASFsNv6JjgBBXYbL+vgnEMc+TxsaWW8ysawQdfpcVocfe2LotYO2JlSCvlyp9f9TuXL
j+S8pTm+ACX5cAxvu5YEFmyBqlHsrSBREsn6CZ6dgUL8kwnkJMaWbNRrl4RsFPK+Aq/yK2y9xRJ+
3JQSSkVinvQnAdjPVtYrIWfa5Lh7pEiNLbhON2ppBoVG+26Z/7JU+WwzpZyASoTvnokY4Grr7cWO
oUF9wOfW0XUx6yNbYV8Gy0we+xKPNPGFyPeL9Cufx1rAIEd57SwI11IvT4HXCG1CLYsxOPTBy5lF
vO977BE2oD/2G7MqvqB7gixt/f0mQo08lvLUq+yVStog21rsI91vgKkr2pJiSf0N3G4aR4hNPHnp
LuqijHfpkGWlnJrX/YXL6gCYHgDpK/DNfy51tGpJIyV2IF+QLjgxdMHmkAhseURcfVo+ULe/g2U6
vdZH4nGIkV0nKZnbzRG14ICrI50l5kDHGpMH1sOGb3RVboFaK8WHAcM0ZAxWepbajhRc4/gdZxg0
lrIrnvCuQgFpFZH6uNsbKJdsMNuENfw+T/S46rvjtPf0EFAAYThK6tNL9FRmZwXftx5wZltxzqxD
eC8wOFgoB1DN8UGOZbu6/PuPLbFQZ7UG1xmnCl+XkosddeRUfLEzKrhNK8o+OELARpr5eHf93OqB
1R1RzUsBWJwjQ1MS1HGv7VZcAadAUVn0Des5VQ6b8eJV+e8tiHTcy1jy8Q7MZ3W1+nWVnWaskC0i
8C917Zit22UVRxiHByMGsSBGxX1tLiHrJTq5NaDwGfFH03N4m24KxKju8WVSEW2XtBeccLuCOSZx
kMjzVwhEyNOPCLmpQVdZZx5qrDG179S3Pz4Gl7vHSgyLmV+PzAxbwlGbmE5NSrZh1GZbAHKCFwTH
zD3TGIyEb0LhvWNeq0+knS8B7XB43OO7BkAzxCX20AlhaOjeMV56Dd7HxCpzOKgNonCj8B9Eh5yC
Ll29LtM3Y1DcIAUlwKX5YcnLws/2CA==
`pragma protect end_protected
